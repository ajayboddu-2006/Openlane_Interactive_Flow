magic
tech sky130A
magscale 1 2
timestamp 1738988163
<< locali >>
rect 9781 13855 9815 14025
<< viali >>
rect 10057 18377 10091 18411
rect 7849 18309 7883 18343
rect 9689 18241 9723 18275
rect 10977 18241 11011 18275
rect 11345 18241 11379 18275
rect 12265 18241 12299 18275
rect 1777 18173 1811 18207
rect 2605 18173 2639 18207
rect 3157 18173 3191 18207
rect 4813 18173 4847 18207
rect 5181 18173 5215 18207
rect 5365 18173 5399 18207
rect 5825 18173 5859 18207
rect 7389 18173 7423 18207
rect 9873 18173 9907 18207
rect 11161 18173 11195 18207
rect 12357 18173 12391 18207
rect 12728 18173 12762 18207
rect 13553 18173 13587 18207
rect 15117 18173 15151 18207
rect 15301 18173 15335 18207
rect 15485 18173 15519 18207
rect 16129 18173 16163 18207
rect 8033 18105 8067 18139
rect 15209 18105 15243 18139
rect 1961 18037 1995 18071
rect 2421 18037 2455 18071
rect 3341 18037 3375 18071
rect 5181 18037 5215 18071
rect 5917 18037 5951 18071
rect 7205 18037 7239 18071
rect 12725 18037 12759 18071
rect 12909 18037 12943 18071
rect 13369 18037 13403 18071
rect 14933 18037 14967 18071
rect 15945 18037 15979 18071
rect 8585 17833 8619 17867
rect 13829 17833 13863 17867
rect 15117 17833 15151 17867
rect 16497 17833 16531 17867
rect 6101 17765 6135 17799
rect 2329 17697 2363 17731
rect 3157 17697 3191 17731
rect 15114 17697 15148 17731
rect 16681 17697 16715 17731
rect 2145 17629 2179 17663
rect 2973 17629 3007 17663
rect 6377 17629 6411 17663
rect 6837 17629 6871 17663
rect 7113 17629 7147 17663
rect 9505 17629 9539 17663
rect 9781 17629 9815 17663
rect 12081 17629 12115 17663
rect 12357 17629 12391 17663
rect 15577 17629 15611 17663
rect 15485 17561 15519 17595
rect 2513 17493 2547 17527
rect 3341 17493 3375 17527
rect 4629 17493 4663 17527
rect 11253 17493 11287 17527
rect 14933 17493 14967 17527
rect 6837 17289 6871 17323
rect 16405 17289 16439 17323
rect 5457 17153 5491 17187
rect 7389 17153 7423 17187
rect 7941 17153 7975 17187
rect 10885 17153 10919 17187
rect 14013 17153 14047 17187
rect 14933 17153 14967 17187
rect 2329 17085 2363 17119
rect 4813 17085 4847 17119
rect 5273 17085 5307 17119
rect 5641 17085 5675 17119
rect 6962 17085 6996 17119
rect 7481 17085 7515 17119
rect 10701 17085 10735 17119
rect 14657 17085 14691 17119
rect 4537 17017 4571 17051
rect 5549 17017 5583 17051
rect 8217 17017 8251 17051
rect 13737 17017 13771 17051
rect 2513 16949 2547 16983
rect 3065 16949 3099 16983
rect 5365 16949 5399 16983
rect 7021 16949 7055 16983
rect 9689 16949 9723 16983
rect 10517 16949 10551 16983
rect 12265 16949 12299 16983
rect 2789 16745 2823 16779
rect 6653 16745 6687 16779
rect 8217 16745 8251 16779
rect 9965 16745 9999 16779
rect 10149 16745 10183 16779
rect 12081 16745 12115 16779
rect 13185 16745 13219 16779
rect 13645 16745 13679 16779
rect 15209 16745 15243 16779
rect 15945 16745 15979 16779
rect 5181 16677 5215 16711
rect 7941 16677 7975 16711
rect 2786 16609 2820 16643
rect 4905 16609 4939 16643
rect 7665 16609 7699 16643
rect 7849 16609 7883 16643
rect 8033 16609 8067 16643
rect 10090 16609 10124 16643
rect 10609 16609 10643 16643
rect 11161 16609 11195 16643
rect 11253 16609 11287 16643
rect 12078 16609 12112 16643
rect 12541 16609 12575 16643
rect 13001 16609 13035 16643
rect 13829 16609 13863 16643
rect 14749 16609 14783 16643
rect 14841 16609 14875 16643
rect 15212 16609 15246 16643
rect 16129 16609 16163 16643
rect 3249 16541 3283 16575
rect 12449 16541 12483 16575
rect 11897 16473 11931 16507
rect 2605 16405 2639 16439
rect 3157 16405 3191 16439
rect 10517 16405 10551 16439
rect 15393 16405 15427 16439
rect 2421 16201 2455 16235
rect 4445 16201 4479 16235
rect 5917 16201 5951 16235
rect 7665 16201 7699 16235
rect 8769 16201 8803 16235
rect 9413 16201 9447 16235
rect 12633 16201 12667 16235
rect 15301 16201 15335 16235
rect 2973 16133 3007 16167
rect 7205 16133 7239 16167
rect 1501 16065 1535 16099
rect 2329 16065 2363 16099
rect 8309 16065 8343 16099
rect 1685 15997 1719 16031
rect 2848 15997 2882 16031
rect 3617 15997 3651 16031
rect 3801 15997 3835 16031
rect 3985 15997 4019 16031
rect 4629 15997 4663 16031
rect 5733 15997 5767 16031
rect 7021 15997 7055 16031
rect 7846 15997 7880 16031
rect 8217 15997 8251 16031
rect 8953 15997 8987 16031
rect 9597 15997 9631 16031
rect 10606 15997 10640 16031
rect 10977 15997 11011 16031
rect 11069 15997 11103 16031
rect 12081 15997 12115 16031
rect 12265 15997 12299 16031
rect 12449 15997 12483 16031
rect 13277 15997 13311 16031
rect 13921 15997 13955 16031
rect 14289 15997 14323 16031
rect 15485 15997 15519 16031
rect 15945 15997 15979 16031
rect 3709 15929 3743 15963
rect 12357 15929 12391 15963
rect 14105 15929 14139 15963
rect 14197 15929 14231 15963
rect 1869 15861 1903 15895
rect 2789 15861 2823 15895
rect 3433 15861 3467 15895
rect 7849 15861 7883 15895
rect 10425 15861 10459 15895
rect 10609 15861 10643 15895
rect 13093 15861 13127 15895
rect 14473 15861 14507 15895
rect 16129 15861 16163 15895
rect 2053 15657 2087 15691
rect 6009 15657 6043 15691
rect 10425 15657 10459 15691
rect 12633 15657 12667 15691
rect 13277 15657 13311 15691
rect 10057 15589 10091 15623
rect 11161 15589 11195 15623
rect 15209 15589 15243 15623
rect 2050 15521 2084 15555
rect 2421 15521 2455 15555
rect 4445 15521 4479 15555
rect 6193 15521 6227 15555
rect 6653 15521 6687 15555
rect 7297 15521 7331 15555
rect 8125 15521 8159 15555
rect 9873 15521 9907 15555
rect 10149 15521 10183 15555
rect 10241 15521 10275 15555
rect 10885 15521 10919 15555
rect 13093 15521 13127 15555
rect 2513 15453 2547 15487
rect 14933 15453 14967 15487
rect 7941 15385 7975 15419
rect 1869 15317 1903 15351
rect 4629 15317 4663 15351
rect 6837 15317 6871 15351
rect 7481 15317 7515 15351
rect 16681 15317 16715 15351
rect 1777 15113 1811 15147
rect 8585 15113 8619 15147
rect 10793 15113 10827 15147
rect 11529 15113 11563 15147
rect 13277 15113 13311 15147
rect 5273 15045 5307 15079
rect 6837 14977 6871 15011
rect 9045 14977 9079 15011
rect 14105 14977 14139 15011
rect 1961 14909 1995 14943
rect 3985 14909 4019 14943
rect 4629 14909 4663 14943
rect 5454 14909 5488 14943
rect 5825 14909 5859 14943
rect 5917 14909 5951 14943
rect 11345 14909 11379 14943
rect 12265 14909 12299 14943
rect 12909 14909 12943 14943
rect 13093 14909 13127 14943
rect 13829 14909 13863 14943
rect 16405 14909 16439 14943
rect 3709 14841 3743 14875
rect 7113 14841 7147 14875
rect 9321 14841 9355 14875
rect 2237 14773 2271 14807
rect 4445 14773 4479 14807
rect 5457 14773 5491 14807
rect 12449 14773 12483 14807
rect 15577 14773 15611 14807
rect 16221 14773 16255 14807
rect 1961 14569 1995 14603
rect 3157 14569 3191 14603
rect 6009 14569 6043 14603
rect 8401 14569 8435 14603
rect 9689 14569 9723 14603
rect 14749 14569 14783 14603
rect 14933 14569 14967 14603
rect 2881 14501 2915 14535
rect 4537 14501 4571 14535
rect 6745 14501 6779 14535
rect 7665 14501 7699 14535
rect 8493 14501 8527 14535
rect 10241 14501 10275 14535
rect 1593 14433 1627 14467
rect 2007 14433 2041 14467
rect 2605 14433 2639 14467
rect 2789 14433 2823 14467
rect 2973 14433 3007 14467
rect 4261 14433 4295 14467
rect 6469 14433 6503 14467
rect 6653 14433 6687 14467
rect 6837 14433 6871 14467
rect 9505 14433 9539 14467
rect 11161 14433 11195 14467
rect 13829 14433 13863 14467
rect 14930 14433 14964 14467
rect 15393 14433 15427 14467
rect 16129 14433 16163 14467
rect 1501 14365 1535 14399
rect 11437 14365 11471 14399
rect 15301 14365 15335 14399
rect 15945 14365 15979 14399
rect 7849 14297 7883 14331
rect 10425 14297 10459 14331
rect 2145 14229 2179 14263
rect 7021 14229 7055 14263
rect 12909 14229 12943 14263
rect 13645 14229 13679 14263
rect 16313 14229 16347 14263
rect 5181 14025 5215 14059
rect 5733 14025 5767 14059
rect 6837 14025 6871 14059
rect 9229 14025 9263 14059
rect 9781 14025 9815 14059
rect 10057 14025 10091 14059
rect 12265 14025 12299 14059
rect 13093 14025 13127 14059
rect 13645 14025 13679 14059
rect 14473 14025 14507 14059
rect 3525 13957 3559 13991
rect 4261 13889 4295 13923
rect 8309 13889 8343 13923
rect 8585 13889 8619 13923
rect 15485 13957 15519 13991
rect 13737 13889 13771 13923
rect 2881 13821 2915 13855
rect 3709 13821 3743 13855
rect 4445 13821 4479 13855
rect 4629 13821 4663 13855
rect 5089 13821 5123 13855
rect 5608 13821 5642 13855
rect 9137 13821 9171 13855
rect 9781 13821 9815 13855
rect 9873 13821 9907 13855
rect 10701 13821 10735 13855
rect 11161 13821 11195 13855
rect 12449 13821 12483 13855
rect 13274 13821 13308 13855
rect 14289 13821 14323 13855
rect 15669 13821 15703 13855
rect 16313 13821 16347 13855
rect 2697 13685 2731 13719
rect 5549 13685 5583 13719
rect 10517 13685 10551 13719
rect 11345 13685 11379 13719
rect 13277 13685 13311 13719
rect 16129 13685 16163 13719
rect 3157 13481 3191 13515
rect 7205 13481 7239 13515
rect 9689 13481 9723 13515
rect 16129 13481 16163 13515
rect 1685 13413 1719 13447
rect 4905 13413 4939 13447
rect 4813 13345 4847 13379
rect 4997 13345 5031 13379
rect 5181 13345 5215 13379
rect 6101 13345 6135 13379
rect 7021 13345 7055 13379
rect 7849 13345 7883 13379
rect 8401 13345 8435 13379
rect 9686 13345 9720 13379
rect 10609 13345 10643 13379
rect 13001 13345 13035 13379
rect 13645 13345 13679 13379
rect 14749 13345 14783 13379
rect 16126 13345 16160 13379
rect 16589 13345 16623 13379
rect 1409 13277 1443 13311
rect 8217 13277 8251 13311
rect 10149 13277 10183 13311
rect 12725 13277 12759 13311
rect 13829 13209 13863 13243
rect 14933 13209 14967 13243
rect 4629 13141 4663 13175
rect 5917 13141 5951 13175
rect 7665 13141 7699 13175
rect 8585 13141 8619 13175
rect 9505 13141 9539 13175
rect 10057 13141 10091 13175
rect 10793 13141 10827 13175
rect 11253 13141 11287 13175
rect 15945 13141 15979 13175
rect 16497 13141 16531 13175
rect 4721 12937 4755 12971
rect 7849 12937 7883 12971
rect 8677 12937 8711 12971
rect 11161 12937 11195 12971
rect 16405 12937 16439 12971
rect 2329 12869 2363 12903
rect 3617 12869 3651 12903
rect 1501 12801 1535 12835
rect 8769 12801 8803 12835
rect 12449 12801 12483 12835
rect 14933 12801 14967 12835
rect 1685 12733 1719 12767
rect 2513 12733 2547 12767
rect 3341 12733 3375 12767
rect 3433 12733 3467 12767
rect 4261 12733 4295 12767
rect 4902 12733 4936 12767
rect 5273 12733 5307 12767
rect 5365 12733 5399 12767
rect 6009 12733 6043 12767
rect 8033 12733 8067 12767
rect 8306 12733 8340 12767
rect 9413 12733 9447 12767
rect 12081 12733 12115 12767
rect 14197 12733 14231 12767
rect 14657 12733 14691 12767
rect 9689 12665 9723 12699
rect 13921 12665 13955 12699
rect 1869 12597 1903 12631
rect 4077 12597 4111 12631
rect 4905 12597 4939 12631
rect 5825 12597 5859 12631
rect 8125 12597 8159 12631
rect 8309 12597 8343 12631
rect 12265 12597 12299 12631
rect 1409 12393 1443 12427
rect 1593 12393 1627 12427
rect 6285 12393 6319 12427
rect 11713 12393 11747 12427
rect 12357 12393 12391 12427
rect 13645 12393 13679 12427
rect 14933 12393 14967 12427
rect 15117 12393 15151 12427
rect 16589 12393 16623 12427
rect 3065 12325 3099 12359
rect 4813 12325 4847 12359
rect 7021 12325 7055 12359
rect 9689 12325 9723 12359
rect 10517 12325 10551 12359
rect 10701 12325 10735 12359
rect 16221 12325 16255 12359
rect 16313 12325 16347 12359
rect 1590 12257 1624 12291
rect 1961 12257 1995 12291
rect 3249 12257 3283 12291
rect 9505 12257 9539 12291
rect 9781 12257 9815 12291
rect 9873 12257 9907 12291
rect 11529 12257 11563 12291
rect 12298 12257 12332 12291
rect 12725 12257 12759 12291
rect 13829 12257 13863 12291
rect 15114 12257 15148 12291
rect 15485 12257 15519 12291
rect 16037 12257 16071 12291
rect 16405 12257 16439 12291
rect 2053 12189 2087 12223
rect 4537 12189 4571 12223
rect 6745 12189 6779 12223
rect 12817 12189 12851 12223
rect 15577 12189 15611 12223
rect 10057 12121 10091 12155
rect 8493 12053 8527 12087
rect 12173 12053 12207 12087
rect 4629 11849 4663 11883
rect 7757 11849 7791 11883
rect 10609 11849 10643 11883
rect 12633 11849 12667 11883
rect 2329 11713 2363 11747
rect 4537 11713 4571 11747
rect 15761 11713 15795 11747
rect 5000 11645 5034 11679
rect 7573 11645 7607 11679
rect 10238 11645 10272 11679
rect 10701 11645 10735 11679
rect 12081 11645 12115 11679
rect 12357 11645 12391 11679
rect 12449 11645 12483 11679
rect 16405 11645 16439 11679
rect 2605 11577 2639 11611
rect 12265 11577 12299 11611
rect 15485 11577 15519 11611
rect 4077 11509 4111 11543
rect 4997 11509 5031 11543
rect 5181 11509 5215 11543
rect 10057 11509 10091 11543
rect 10241 11509 10275 11543
rect 14013 11509 14047 11543
rect 16221 11509 16255 11543
rect 2145 11305 2179 11339
rect 2329 11305 2363 11339
rect 6285 11305 6319 11339
rect 7113 11305 7147 11339
rect 12265 11305 12299 11339
rect 13829 11305 13863 11339
rect 16681 11305 16715 11339
rect 4813 11237 4847 11271
rect 1777 11169 1811 11203
rect 2326 11169 2360 11203
rect 2789 11169 2823 11203
rect 7110 11169 7144 11203
rect 8585 11169 8619 11203
rect 11897 11169 11931 11203
rect 12268 11169 12302 11203
rect 12909 11169 12943 11203
rect 13645 11169 13679 11203
rect 14933 11169 14967 11203
rect 4537 11101 4571 11135
rect 7573 11101 7607 11135
rect 9597 11101 9631 11135
rect 11069 11101 11103 11135
rect 11345 11101 11379 11135
rect 11805 11101 11839 11135
rect 1961 11033 1995 11067
rect 7481 11033 7515 11067
rect 8401 11033 8435 11067
rect 13093 11033 13127 11067
rect 2697 10965 2731 10999
rect 6929 10965 6963 10999
rect 12449 10965 12483 10999
rect 15196 10965 15230 10999
rect 2605 10761 2639 10795
rect 5457 10761 5491 10795
rect 10149 10761 10183 10795
rect 10885 10761 10919 10795
rect 11345 10761 11379 10795
rect 15393 10761 15427 10795
rect 9597 10693 9631 10727
rect 3709 10625 3743 10659
rect 3985 10625 4019 10659
rect 12081 10625 12115 10659
rect 12357 10625 12391 10659
rect 13829 10625 13863 10659
rect 14381 10625 14415 10659
rect 2053 10557 2087 10591
rect 2237 10557 2271 10591
rect 2421 10557 2455 10591
rect 3249 10557 3283 10591
rect 9137 10557 9171 10591
rect 9722 10557 9756 10591
rect 10241 10557 10275 10591
rect 10333 10557 10367 10591
rect 10517 10557 10551 10591
rect 10701 10557 10735 10591
rect 11529 10557 11563 10591
rect 14289 10557 14323 10591
rect 14752 10557 14786 10591
rect 15577 10557 15611 10591
rect 15669 10557 15703 10591
rect 15761 10557 15795 10591
rect 15945 10557 15979 10591
rect 2329 10489 2363 10523
rect 8861 10489 8895 10523
rect 10609 10489 10643 10523
rect 3065 10421 3099 10455
rect 7389 10421 7423 10455
rect 9781 10421 9815 10455
rect 14749 10421 14783 10455
rect 14933 10421 14967 10455
rect 3157 10217 3191 10251
rect 5181 10217 5215 10251
rect 5825 10217 5859 10251
rect 6837 10217 6871 10251
rect 7021 10217 7055 10251
rect 8493 10217 8527 10251
rect 11713 10217 11747 10251
rect 13185 10217 13219 10251
rect 1685 10149 1719 10183
rect 8217 10149 8251 10183
rect 15669 10149 15703 10183
rect 5365 10081 5399 10115
rect 6009 10081 6043 10115
rect 7018 10081 7052 10115
rect 7941 10081 7975 10115
rect 8125 10081 8159 10115
rect 8309 10081 8343 10115
rect 9505 10081 9539 10115
rect 11897 10081 11931 10115
rect 12081 10081 12115 10115
rect 13182 10081 13216 10115
rect 13553 10081 13587 10115
rect 15485 10081 15519 10115
rect 15577 10081 15611 10115
rect 15853 10081 15887 10115
rect 16497 10081 16531 10115
rect 1409 10013 1443 10047
rect 7389 10013 7423 10047
rect 7481 10013 7515 10047
rect 13645 10013 13679 10047
rect 10793 9945 10827 9979
rect 13001 9877 13035 9911
rect 15301 9877 15335 9911
rect 16313 9877 16347 9911
rect 5917 9673 5951 9707
rect 15853 9673 15887 9707
rect 7389 9605 7423 9639
rect 9965 9537 9999 9571
rect 10977 9537 11011 9571
rect 11069 9537 11103 9571
rect 13001 9537 13035 9571
rect 13277 9537 13311 9571
rect 14749 9537 14783 9571
rect 15301 9537 15335 9571
rect 3617 9469 3651 9503
rect 4629 9469 4663 9503
rect 5273 9469 5307 9503
rect 5365 9469 5399 9503
rect 5736 9469 5770 9503
rect 7018 9469 7052 9503
rect 7481 9469 7515 9503
rect 8217 9469 8251 9503
rect 10606 9469 10640 9503
rect 12265 9469 12299 9503
rect 15209 9469 15243 9503
rect 15728 9469 15762 9503
rect 8493 9401 8527 9435
rect 3801 9333 3835 9367
rect 4813 9333 4847 9367
rect 5733 9333 5767 9367
rect 6837 9333 6871 9367
rect 7021 9333 7055 9367
rect 10425 9333 10459 9367
rect 10609 9333 10643 9367
rect 12081 9333 12115 9367
rect 15669 9333 15703 9367
rect 1409 9129 1443 9163
rect 1593 9129 1627 9163
rect 2697 9129 2731 9163
rect 8217 9129 8251 9163
rect 12357 9129 12391 9163
rect 13185 9129 13219 9163
rect 13829 9129 13863 9163
rect 16681 9129 16715 9163
rect 9873 9061 9907 9095
rect 15209 9061 15243 9095
rect 1590 8993 1624 9027
rect 2694 8993 2728 9027
rect 3157 8993 3191 9027
rect 9597 8993 9631 9027
rect 9781 8993 9815 9027
rect 9965 8993 9999 9027
rect 13001 8993 13035 9027
rect 13645 8993 13679 9027
rect 14933 8993 14967 9027
rect 2053 8925 2087 8959
rect 5733 8925 5767 8959
rect 6009 8925 6043 8959
rect 6469 8925 6503 8959
rect 6745 8925 6779 8959
rect 10609 8925 10643 8959
rect 10885 8925 10919 8959
rect 12817 8925 12851 8959
rect 10149 8857 10183 8891
rect 1961 8789 1995 8823
rect 2513 8789 2547 8823
rect 3065 8789 3099 8823
rect 4261 8789 4295 8823
rect 2605 8585 2639 8619
rect 7389 8585 7423 8619
rect 7849 8585 7883 8619
rect 9045 8585 9079 8619
rect 10425 8585 10459 8619
rect 10977 8585 11011 8619
rect 12265 8585 12299 8619
rect 15117 8585 15151 8619
rect 15669 8585 15703 8619
rect 4997 8517 5031 8551
rect 1869 8449 1903 8483
rect 4353 8449 4387 8483
rect 14289 8449 14323 8483
rect 14565 8449 14599 8483
rect 1685 8381 1719 8415
rect 4813 8381 4847 8415
rect 5641 8381 5675 8415
rect 6101 8381 6135 8415
rect 6837 8381 6871 8415
rect 7113 8381 7147 8415
rect 7205 8381 7239 8415
rect 8033 8381 8067 8415
rect 8125 8381 8159 8415
rect 8677 8381 8711 8415
rect 8861 8381 8895 8415
rect 10026 8381 10060 8415
rect 10517 8381 10551 8415
rect 11161 8381 11195 8415
rect 12081 8381 12115 8415
rect 15270 8381 15304 8415
rect 15761 8381 15795 8415
rect 16405 8381 16439 8415
rect 4077 8313 4111 8347
rect 7021 8313 7055 8347
rect 10122 8313 10156 8347
rect 15366 8313 15400 8347
rect 1501 8245 1535 8279
rect 5457 8245 5491 8279
rect 6285 8245 6319 8279
rect 9873 8245 9907 8279
rect 12817 8245 12851 8279
rect 16221 8245 16255 8279
rect 1777 8041 1811 8075
rect 2881 8041 2915 8075
rect 5457 8041 5491 8075
rect 11529 8041 11563 8075
rect 12173 8041 12207 8075
rect 13829 8041 13863 8075
rect 14933 8041 14967 8075
rect 15577 8041 15611 8075
rect 2605 7973 2639 8007
rect 8033 7973 8067 8007
rect 8217 7973 8251 8007
rect 10057 7973 10091 8007
rect 1961 7905 1995 7939
rect 2329 7905 2363 7939
rect 2513 7905 2547 7939
rect 2697 7905 2731 7939
rect 4445 7905 4479 7939
rect 4537 7905 4571 7939
rect 5273 7905 5307 7939
rect 9505 7905 9539 7939
rect 12170 7905 12204 7939
rect 13645 7905 13679 7939
rect 14749 7905 14783 7939
rect 15761 7905 15795 7939
rect 15853 7905 15887 7939
rect 16681 7905 16715 7939
rect 5089 7837 5123 7871
rect 9781 7837 9815 7871
rect 12633 7837 12667 7871
rect 16497 7769 16531 7803
rect 4261 7701 4295 7735
rect 9689 7701 9723 7735
rect 11989 7701 12023 7735
rect 12541 7701 12575 7735
rect 2605 7497 2639 7531
rect 3709 7497 3743 7531
rect 10517 7497 10551 7531
rect 10977 7497 11011 7531
rect 15669 7497 15703 7531
rect 3157 7429 3191 7463
rect 7481 7429 7515 7463
rect 7849 7429 7883 7463
rect 8953 7429 8987 7463
rect 2697 7361 2731 7395
rect 5917 7361 5951 7395
rect 7757 7361 7791 7395
rect 10149 7361 10183 7395
rect 12081 7361 12115 7395
rect 2234 7293 2268 7327
rect 3282 7293 3316 7327
rect 3801 7293 3835 7327
rect 4445 7293 4479 7327
rect 4629 7293 4663 7327
rect 4813 7293 4847 7327
rect 5454 7293 5488 7327
rect 5825 7293 5859 7327
rect 7021 7293 7055 7327
rect 7665 7293 7699 7327
rect 8220 7293 8254 7327
rect 8861 7293 8895 7327
rect 9380 7293 9414 7327
rect 10333 7293 10367 7327
rect 11161 7293 11195 7327
rect 12265 7293 12299 7327
rect 13001 7293 13035 7327
rect 15853 7293 15887 7327
rect 15945 7293 15979 7327
rect 4537 7225 4571 7259
rect 13277 7225 13311 7259
rect 2053 7157 2087 7191
rect 2237 7157 2271 7191
rect 3341 7157 3375 7191
rect 4261 7157 4295 7191
rect 5273 7157 5307 7191
rect 5457 7157 5491 7191
rect 6837 7157 6871 7191
rect 8217 7157 8251 7191
rect 8401 7157 8435 7191
rect 9321 7157 9355 7191
rect 9505 7157 9539 7191
rect 12449 7157 12483 7191
rect 14749 7157 14783 7191
rect 12357 6953 12391 6987
rect 12541 6953 12575 6987
rect 1685 6885 1719 6919
rect 4813 6885 4847 6919
rect 13185 6885 13219 6919
rect 6745 6817 6779 6851
rect 9505 6817 9539 6851
rect 10333 6817 10367 6851
rect 10793 6817 10827 6851
rect 11897 6817 11931 6851
rect 12360 6817 12394 6851
rect 13001 6817 13035 6851
rect 13277 6817 13311 6851
rect 13369 6817 13403 6851
rect 15117 6817 15151 6851
rect 15301 6817 15335 6851
rect 15393 6817 15427 6851
rect 15531 6817 15565 6851
rect 16313 6817 16347 6851
rect 1409 6749 1443 6783
rect 3157 6749 3191 6783
rect 4537 6749 4571 6783
rect 7021 6749 7055 6783
rect 8493 6749 8527 6783
rect 11989 6749 12023 6783
rect 16497 6749 16531 6783
rect 10149 6681 10183 6715
rect 13553 6681 13587 6715
rect 16129 6681 16163 6715
rect 6285 6613 6319 6647
rect 9689 6613 9723 6647
rect 10977 6613 11011 6647
rect 15669 6613 15703 6647
rect 2421 6409 2455 6443
rect 3157 6409 3191 6443
rect 7941 6409 7975 6443
rect 13369 6409 13403 6443
rect 13921 6409 13955 6443
rect 14933 6409 14967 6443
rect 15485 6409 15519 6443
rect 16221 6409 16255 6443
rect 4629 6273 4663 6307
rect 9321 6273 9355 6307
rect 2237 6205 2271 6239
rect 4905 6205 4939 6239
rect 5365 6205 5399 6239
rect 5549 6205 5583 6239
rect 7113 6205 7147 6239
rect 8125 6205 8159 6239
rect 8217 6205 8251 6239
rect 8493 6205 8527 6239
rect 9045 6205 9079 6239
rect 12081 6205 12115 6239
rect 13185 6205 13219 6239
rect 13829 6205 13863 6239
rect 14348 6205 14382 6239
rect 15114 6205 15148 6239
rect 15577 6205 15611 6239
rect 16405 6205 16439 6239
rect 8309 6137 8343 6171
rect 5733 6069 5767 6103
rect 6929 6069 6963 6103
rect 10793 6069 10827 6103
rect 12265 6069 12299 6103
rect 14289 6069 14323 6103
rect 14473 6069 14507 6103
rect 15117 6069 15151 6103
rect 1593 5865 1627 5899
rect 4261 5865 4295 5899
rect 5641 5865 5675 5899
rect 10701 5865 10735 5899
rect 11529 5865 11563 5899
rect 13829 5865 13863 5899
rect 16681 5865 16715 5899
rect 8309 5797 8343 5831
rect 15209 5797 15243 5831
rect 1409 5729 1443 5763
rect 4445 5729 4479 5763
rect 5825 5729 5859 5763
rect 10057 5729 10091 5763
rect 10885 5729 10919 5763
rect 11526 5729 11560 5763
rect 12587 5729 12621 5763
rect 12725 5729 12759 5763
rect 12817 5729 12851 5763
rect 13001 5729 13035 5763
rect 13645 5729 13679 5763
rect 7389 5661 7423 5695
rect 7665 5661 7699 5695
rect 9873 5661 9907 5695
rect 11897 5661 11931 5695
rect 11989 5661 12023 5695
rect 14933 5661 14967 5695
rect 11345 5593 11379 5627
rect 5917 5525 5951 5559
rect 8217 5525 8251 5559
rect 10241 5525 10275 5559
rect 12449 5525 12483 5559
rect 3709 5321 3743 5355
rect 4353 5321 4387 5355
rect 5273 5321 5307 5355
rect 6837 5321 6871 5355
rect 11069 5321 11103 5355
rect 13829 5321 13863 5355
rect 5825 5185 5859 5219
rect 12081 5185 12115 5219
rect 12357 5185 12391 5219
rect 14289 5185 14323 5219
rect 14565 5185 14599 5219
rect 1961 5117 1995 5151
rect 4169 5117 4203 5151
rect 5454 5117 5488 5151
rect 5917 5117 5951 5151
rect 7021 5117 7055 5151
rect 7205 5117 7239 5151
rect 7389 5117 7423 5151
rect 7941 5117 7975 5151
rect 10698 5117 10732 5151
rect 11161 5117 11195 5151
rect 2237 5049 2271 5083
rect 7113 5049 7147 5083
rect 8217 5049 8251 5083
rect 5457 4981 5491 5015
rect 9689 4981 9723 5015
rect 10517 4981 10551 5015
rect 10701 4981 10735 5015
rect 16037 4981 16071 5015
rect 2973 4777 3007 4811
rect 6009 4777 6043 4811
rect 9505 4777 9539 4811
rect 12817 4777 12851 4811
rect 13277 4777 13311 4811
rect 14933 4777 14967 4811
rect 16221 4777 16255 4811
rect 10517 4709 10551 4743
rect 2789 4641 2823 4675
rect 4261 4641 4295 4675
rect 7205 4641 7239 4675
rect 8585 4641 8619 4675
rect 9689 4641 9723 4675
rect 10241 4641 10275 4675
rect 12633 4641 12667 4675
rect 13461 4641 13495 4675
rect 14749 4641 14783 4675
rect 15761 4641 15795 4675
rect 16405 4641 16439 4675
rect 4537 4573 4571 4607
rect 8309 4573 8343 4607
rect 12449 4573 12483 4607
rect 7021 4437 7055 4471
rect 11989 4437 12023 4471
rect 15577 4437 15611 4471
rect 5641 4233 5675 4267
rect 8033 4233 8067 4267
rect 10977 4233 11011 4267
rect 12081 4233 12115 4267
rect 15669 4233 15703 4267
rect 6837 4165 6871 4199
rect 8677 4165 8711 4199
rect 9321 4097 9355 4131
rect 14473 4097 14507 4131
rect 3249 4029 3283 4063
rect 3893 4029 3927 4063
rect 4997 4029 5031 4063
rect 5181 4029 5215 4063
rect 5825 4029 5859 4063
rect 7021 4029 7055 4063
rect 8125 4029 8159 4063
rect 8861 4029 8895 4063
rect 9413 4029 9447 4063
rect 9784 4029 9818 4063
rect 10425 4029 10459 4063
rect 10609 4029 10643 4063
rect 10701 4029 10735 4063
rect 10793 4029 10827 4063
rect 12265 4029 12299 4063
rect 15298 4029 15332 4063
rect 15761 4029 15795 4063
rect 16397 4029 16431 4063
rect 14197 3961 14231 3995
rect 3433 3893 3467 3927
rect 4077 3893 4111 3927
rect 4813 3893 4847 3927
rect 9781 3893 9815 3927
rect 9965 3893 9999 3927
rect 12725 3893 12759 3927
rect 15117 3893 15151 3927
rect 15301 3893 15335 3927
rect 16221 3893 16255 3927
rect 2697 3689 2731 3723
rect 2881 3689 2915 3723
rect 4813 3689 4847 3723
rect 4997 3689 5031 3723
rect 9689 3689 9723 3723
rect 10793 3689 10827 3723
rect 13737 3689 13771 3723
rect 2053 3553 2087 3587
rect 2878 3553 2912 3587
rect 4994 3553 5028 3587
rect 8401 3553 8435 3587
rect 9686 3553 9720 3587
rect 10057 3553 10091 3587
rect 10149 3553 10183 3587
rect 10609 3553 10643 3587
rect 11437 3553 11471 3587
rect 11621 3553 11655 3587
rect 11713 3553 11747 3587
rect 11851 3553 11885 3587
rect 12633 3553 12667 3587
rect 13553 3553 13587 3587
rect 14933 3553 14967 3587
rect 3249 3485 3283 3519
rect 3341 3485 3375 3519
rect 5457 3485 5491 3519
rect 7389 3485 7423 3519
rect 7665 3485 7699 3519
rect 15209 3485 15243 3519
rect 16681 3485 16715 3519
rect 11989 3417 12023 3451
rect 2237 3349 2271 3383
rect 5365 3349 5399 3383
rect 5917 3349 5951 3383
rect 8217 3349 8251 3383
rect 9505 3349 9539 3383
rect 12449 3349 12483 3383
rect 1961 3145 1995 3179
rect 4537 3145 4571 3179
rect 9229 3145 9263 3179
rect 12081 3145 12115 3179
rect 13829 3145 13863 3179
rect 14473 3145 14507 3179
rect 15025 3145 15059 3179
rect 16129 3145 16163 3179
rect 2329 3009 2363 3043
rect 4077 3009 4111 3043
rect 5089 3009 5123 3043
rect 7021 3009 7055 3043
rect 8493 3009 8527 3043
rect 8769 3009 8803 3043
rect 10977 3009 11011 3043
rect 12725 3009 12759 3043
rect 1777 2941 1811 2975
rect 4662 2941 4696 2975
rect 5181 2941 5215 2975
rect 12262 2941 12296 2975
rect 12633 2941 12667 2975
rect 13369 2941 13403 2975
rect 14013 2941 14047 2975
rect 14654 2941 14688 2975
rect 15117 2941 15151 2975
rect 15577 2941 15611 2975
rect 15853 2941 15887 2975
rect 15945 2941 15979 2975
rect 2605 2873 2639 2907
rect 5733 2873 5767 2907
rect 10701 2873 10735 2907
rect 15761 2873 15795 2907
rect 4721 2805 4755 2839
rect 5825 2805 5859 2839
rect 12265 2805 12299 2839
rect 13185 2805 13219 2839
rect 14657 2805 14691 2839
rect 2973 2601 3007 2635
rect 4813 2601 4847 2635
rect 5549 2601 5583 2635
rect 7481 2601 7515 2635
rect 8677 2601 8711 2635
rect 10517 2601 10551 2635
rect 10701 2601 10735 2635
rect 12265 2601 12299 2635
rect 15485 2601 15519 2635
rect 4537 2533 4571 2567
rect 7113 2533 7147 2567
rect 7205 2533 7239 2567
rect 13737 2533 13771 2567
rect 1961 2465 1995 2499
rect 3157 2465 3191 2499
rect 4261 2465 4295 2499
rect 4445 2465 4479 2499
rect 4629 2465 4663 2499
rect 5546 2465 5580 2499
rect 6009 2465 6043 2499
rect 6929 2465 6963 2499
rect 7297 2465 7331 2499
rect 8493 2465 8527 2499
rect 9781 2465 9815 2499
rect 9873 2465 9907 2499
rect 10057 2465 10091 2499
rect 10698 2465 10732 2499
rect 11161 2465 11195 2499
rect 14013 2465 14047 2499
rect 15669 2465 15703 2499
rect 15761 2465 15795 2499
rect 16681 2465 16715 2499
rect 3341 2397 3375 2431
rect 2145 2329 2179 2363
rect 5365 2329 5399 2363
rect 11069 2329 11103 2363
rect 5917 2261 5951 2295
rect 16497 2261 16531 2295
<< metal1 >>
rect 1104 18522 17388 18544
rect 1104 18470 3696 18522
rect 3748 18470 3760 18522
rect 3812 18470 3824 18522
rect 3876 18470 3888 18522
rect 3940 18470 9124 18522
rect 9176 18470 9188 18522
rect 9240 18470 9252 18522
rect 9304 18470 9316 18522
rect 9368 18470 14552 18522
rect 14604 18470 14616 18522
rect 14668 18470 14680 18522
rect 14732 18470 14744 18522
rect 14796 18470 17388 18522
rect 1104 18448 17388 18470
rect 10045 18411 10103 18417
rect 10045 18377 10057 18411
rect 10091 18408 10103 18411
rect 15286 18408 15292 18420
rect 10091 18380 15292 18408
rect 10091 18377 10103 18380
rect 10045 18371 10103 18377
rect 15286 18368 15292 18380
rect 15344 18368 15350 18420
rect 7834 18340 7840 18352
rect 7795 18312 7840 18340
rect 7834 18300 7840 18312
rect 7892 18300 7898 18352
rect 16482 18340 16488 18352
rect 11164 18312 16488 18340
rect 934 18232 940 18284
rect 992 18272 998 18284
rect 9677 18275 9735 18281
rect 992 18244 2636 18272
rect 992 18232 998 18244
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 2608 18213 2636 18244
rect 9677 18241 9689 18275
rect 9723 18272 9735 18275
rect 10134 18272 10140 18284
rect 9723 18244 10140 18272
rect 9723 18241 9735 18244
rect 9677 18235 9735 18241
rect 10134 18232 10140 18244
rect 10192 18272 10198 18284
rect 10965 18275 11023 18281
rect 10965 18272 10977 18275
rect 10192 18244 10977 18272
rect 10192 18232 10198 18244
rect 10965 18241 10977 18244
rect 11011 18241 11023 18275
rect 10965 18235 11023 18241
rect 2593 18207 2651 18213
rect 2593 18173 2605 18207
rect 2639 18173 2651 18207
rect 2593 18167 2651 18173
rect 3145 18207 3203 18213
rect 3145 18173 3157 18207
rect 3191 18204 3203 18207
rect 4062 18204 4068 18216
rect 3191 18176 4068 18204
rect 3191 18173 3203 18176
rect 3145 18167 3203 18173
rect 4062 18164 4068 18176
rect 4120 18164 4126 18216
rect 4798 18204 4804 18216
rect 4759 18176 4804 18204
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 5074 18164 5080 18216
rect 5132 18204 5138 18216
rect 5169 18207 5227 18213
rect 5169 18204 5181 18207
rect 5132 18176 5181 18204
rect 5132 18164 5138 18176
rect 5169 18173 5181 18176
rect 5215 18173 5227 18207
rect 5169 18167 5227 18173
rect 5353 18207 5411 18213
rect 5353 18173 5365 18207
rect 5399 18204 5411 18207
rect 5534 18204 5540 18216
rect 5399 18176 5540 18204
rect 5399 18173 5411 18176
rect 5353 18167 5411 18173
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 5813 18207 5871 18213
rect 5813 18173 5825 18207
rect 5859 18173 5871 18207
rect 5813 18167 5871 18173
rect 7377 18207 7435 18213
rect 7377 18173 7389 18207
rect 7423 18204 7435 18207
rect 8938 18204 8944 18216
rect 7423 18176 8944 18204
rect 7423 18173 7435 18176
rect 7377 18167 7435 18173
rect 5258 18136 5264 18148
rect 5171 18108 5264 18136
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 2314 18028 2320 18080
rect 2372 18068 2378 18080
rect 2409 18071 2467 18077
rect 2409 18068 2421 18071
rect 2372 18040 2421 18068
rect 2372 18028 2378 18040
rect 2409 18037 2421 18040
rect 2455 18037 2467 18071
rect 2409 18031 2467 18037
rect 3329 18071 3387 18077
rect 3329 18037 3341 18071
rect 3375 18068 3387 18071
rect 4706 18068 4712 18080
rect 3375 18040 4712 18068
rect 3375 18037 3387 18040
rect 3329 18031 3387 18037
rect 4706 18028 4712 18040
rect 4764 18028 4770 18080
rect 5184 18077 5212 18108
rect 5258 18096 5264 18108
rect 5316 18136 5322 18148
rect 5828 18136 5856 18167
rect 8938 18164 8944 18176
rect 8996 18164 9002 18216
rect 9858 18204 9864 18216
rect 9819 18176 9864 18204
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 11164 18213 11192 18312
rect 16482 18300 16488 18312
rect 16540 18300 16546 18352
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18272 11391 18275
rect 12158 18272 12164 18284
rect 11379 18244 12164 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 12158 18232 12164 18244
rect 12216 18272 12222 18284
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 12216 18244 12265 18272
rect 12216 18232 12222 18244
rect 12253 18241 12265 18244
rect 12299 18272 12311 18275
rect 12299 18244 12480 18272
rect 12299 18241 12311 18244
rect 12253 18235 12311 18241
rect 11149 18207 11207 18213
rect 11149 18173 11161 18207
rect 11195 18173 11207 18207
rect 12342 18204 12348 18216
rect 12303 18176 12348 18204
rect 11149 18167 11207 18173
rect 12342 18164 12348 18176
rect 12400 18164 12406 18216
rect 12452 18204 12480 18244
rect 12894 18232 12900 18284
rect 12952 18272 12958 18284
rect 12952 18244 16160 18272
rect 12952 18232 12958 18244
rect 12716 18207 12774 18213
rect 12716 18204 12728 18207
rect 12452 18176 12728 18204
rect 12716 18173 12728 18176
rect 12762 18173 12774 18207
rect 12716 18167 12774 18173
rect 13541 18207 13599 18213
rect 13541 18173 13553 18207
rect 13587 18173 13599 18207
rect 15102 18204 15108 18216
rect 15063 18176 15108 18204
rect 13541 18167 13599 18173
rect 5316 18108 5856 18136
rect 8021 18139 8079 18145
rect 5316 18096 5322 18108
rect 8021 18105 8033 18139
rect 8067 18136 8079 18139
rect 8570 18136 8576 18148
rect 8067 18108 8576 18136
rect 8067 18105 8079 18108
rect 8021 18099 8079 18105
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 11054 18096 11060 18148
rect 11112 18136 11118 18148
rect 13556 18136 13584 18167
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 15286 18204 15292 18216
rect 15247 18176 15292 18204
rect 15286 18164 15292 18176
rect 15344 18164 15350 18216
rect 15378 18164 15384 18216
rect 15436 18204 15442 18216
rect 16132 18213 16160 18244
rect 15473 18207 15531 18213
rect 15473 18204 15485 18207
rect 15436 18176 15485 18204
rect 15436 18164 15442 18176
rect 15473 18173 15485 18176
rect 15519 18173 15531 18207
rect 15473 18167 15531 18173
rect 16117 18207 16175 18213
rect 16117 18173 16129 18207
rect 16163 18173 16175 18207
rect 16117 18167 16175 18173
rect 15194 18136 15200 18148
rect 11112 18108 13584 18136
rect 15155 18108 15200 18136
rect 11112 18096 11118 18108
rect 15194 18096 15200 18108
rect 15252 18096 15258 18148
rect 5169 18071 5227 18077
rect 5169 18037 5181 18071
rect 5215 18037 5227 18071
rect 5169 18031 5227 18037
rect 5905 18071 5963 18077
rect 5905 18037 5917 18071
rect 5951 18068 5963 18071
rect 6086 18068 6092 18080
rect 5951 18040 6092 18068
rect 5951 18037 5963 18040
rect 5905 18031 5963 18037
rect 6086 18028 6092 18040
rect 6144 18028 6150 18080
rect 6822 18028 6828 18080
rect 6880 18068 6886 18080
rect 7193 18071 7251 18077
rect 7193 18068 7205 18071
rect 6880 18040 7205 18068
rect 6880 18028 6886 18040
rect 7193 18037 7205 18040
rect 7239 18037 7251 18071
rect 7193 18031 7251 18037
rect 12342 18028 12348 18080
rect 12400 18068 12406 18080
rect 12713 18071 12771 18077
rect 12713 18068 12725 18071
rect 12400 18040 12725 18068
rect 12400 18028 12406 18040
rect 12713 18037 12725 18040
rect 12759 18037 12771 18071
rect 12894 18068 12900 18080
rect 12855 18040 12900 18068
rect 12713 18031 12771 18037
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 13354 18068 13360 18080
rect 13315 18040 13360 18068
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 14918 18068 14924 18080
rect 14879 18040 14924 18068
rect 14918 18028 14924 18040
rect 14976 18028 14982 18080
rect 15470 18028 15476 18080
rect 15528 18068 15534 18080
rect 15933 18071 15991 18077
rect 15933 18068 15945 18071
rect 15528 18040 15945 18068
rect 15528 18028 15534 18040
rect 15933 18037 15945 18040
rect 15979 18037 15991 18071
rect 15933 18031 15991 18037
rect 1104 17978 17388 18000
rect 1104 17926 6410 17978
rect 6462 17926 6474 17978
rect 6526 17926 6538 17978
rect 6590 17926 6602 17978
rect 6654 17926 11838 17978
rect 11890 17926 11902 17978
rect 11954 17926 11966 17978
rect 12018 17926 12030 17978
rect 12082 17926 17388 17978
rect 1104 17904 17388 17926
rect 6822 17864 6828 17876
rect 5644 17836 6828 17864
rect 1946 17756 1952 17808
rect 2004 17796 2010 17808
rect 2004 17768 2774 17796
rect 5644 17782 5672 17836
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 8570 17864 8576 17876
rect 8531 17836 8576 17864
rect 8570 17824 8576 17836
rect 8628 17824 8634 17876
rect 13817 17867 13875 17873
rect 13817 17833 13829 17867
rect 13863 17864 13875 17867
rect 15102 17864 15108 17876
rect 13863 17836 15108 17864
rect 13863 17833 13875 17836
rect 13817 17827 13875 17833
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 16482 17864 16488 17876
rect 16443 17836 16488 17864
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 6086 17796 6092 17808
rect 6047 17768 6092 17796
rect 2004 17756 2010 17768
rect 2314 17728 2320 17740
rect 2275 17700 2320 17728
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 2746 17728 2774 17768
rect 6086 17756 6092 17768
rect 6144 17756 6150 17808
rect 8754 17796 8760 17808
rect 8326 17768 8760 17796
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 10042 17756 10048 17808
rect 10100 17796 10106 17808
rect 13630 17796 13636 17808
rect 10100 17768 10258 17796
rect 13570 17768 13636 17796
rect 10100 17756 10106 17768
rect 13630 17756 13636 17768
rect 13688 17756 13694 17808
rect 3145 17731 3203 17737
rect 3145 17728 3157 17731
rect 2746 17700 3157 17728
rect 3145 17697 3157 17700
rect 3191 17697 3203 17731
rect 3145 17691 3203 17697
rect 15102 17731 15160 17737
rect 15102 17697 15114 17731
rect 15148 17728 15160 17731
rect 15194 17728 15200 17740
rect 15148 17700 15200 17728
rect 15148 17697 15160 17700
rect 15102 17691 15160 17697
rect 15194 17688 15200 17700
rect 15252 17728 15258 17740
rect 16669 17731 16727 17737
rect 15252 17700 15608 17728
rect 15252 17688 15258 17700
rect 15580 17672 15608 17700
rect 16669 17697 16681 17731
rect 16715 17728 16727 17731
rect 17954 17728 17960 17740
rect 16715 17700 17960 17728
rect 16715 17697 16727 17700
rect 16669 17691 16727 17697
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17660 2191 17663
rect 2961 17663 3019 17669
rect 2961 17660 2973 17663
rect 2179 17632 2973 17660
rect 2179 17629 2191 17632
rect 2133 17623 2191 17629
rect 2961 17629 2973 17632
rect 3007 17660 3019 17663
rect 3510 17660 3516 17672
rect 3007 17632 3516 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 3510 17620 3516 17632
rect 3568 17660 3574 17672
rect 5074 17660 5080 17672
rect 3568 17632 5080 17660
rect 3568 17620 3574 17632
rect 5074 17620 5080 17632
rect 5132 17620 5138 17672
rect 6365 17663 6423 17669
rect 6365 17629 6377 17663
rect 6411 17660 6423 17663
rect 6730 17660 6736 17672
rect 6411 17632 6736 17660
rect 6411 17629 6423 17632
rect 6365 17623 6423 17629
rect 6730 17620 6736 17632
rect 6788 17660 6794 17672
rect 6825 17663 6883 17669
rect 6825 17660 6837 17663
rect 6788 17632 6837 17660
rect 6788 17620 6794 17632
rect 6825 17629 6837 17632
rect 6871 17629 6883 17663
rect 7098 17660 7104 17672
rect 7059 17632 7104 17660
rect 6825 17623 6883 17629
rect 7098 17620 7104 17632
rect 7156 17620 7162 17672
rect 9493 17663 9551 17669
rect 9493 17629 9505 17663
rect 9539 17660 9551 17663
rect 9766 17660 9772 17672
rect 9539 17632 9628 17660
rect 9727 17632 9772 17660
rect 9539 17629 9551 17632
rect 9493 17623 9551 17629
rect 2498 17524 2504 17536
rect 2459 17496 2504 17524
rect 2498 17484 2504 17496
rect 2556 17484 2562 17536
rect 3326 17524 3332 17536
rect 3287 17496 3332 17524
rect 3326 17484 3332 17496
rect 3384 17484 3390 17536
rect 4617 17527 4675 17533
rect 4617 17493 4629 17527
rect 4663 17524 4675 17527
rect 4798 17524 4804 17536
rect 4663 17496 4804 17524
rect 4663 17493 4675 17496
rect 4617 17487 4675 17493
rect 4798 17484 4804 17496
rect 4856 17524 4862 17536
rect 5350 17524 5356 17536
rect 4856 17496 5356 17524
rect 4856 17484 4862 17496
rect 5350 17484 5356 17496
rect 5408 17484 5414 17536
rect 9600 17524 9628 17632
rect 9766 17620 9772 17632
rect 9824 17620 9830 17672
rect 12069 17663 12127 17669
rect 12069 17660 12081 17663
rect 10796 17632 12081 17660
rect 10796 17524 10824 17632
rect 12069 17629 12081 17632
rect 12115 17629 12127 17663
rect 12069 17623 12127 17629
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17660 12403 17663
rect 12894 17660 12900 17672
rect 12391 17632 12900 17660
rect 12391 17629 12403 17632
rect 12345 17623 12403 17629
rect 12894 17620 12900 17632
rect 12952 17620 12958 17672
rect 15562 17660 15568 17672
rect 15523 17632 15568 17660
rect 15562 17620 15568 17632
rect 15620 17620 15626 17672
rect 15102 17552 15108 17604
rect 15160 17592 15166 17604
rect 15473 17595 15531 17601
rect 15473 17592 15485 17595
rect 15160 17564 15485 17592
rect 15160 17552 15166 17564
rect 15473 17561 15485 17564
rect 15519 17561 15531 17595
rect 15473 17555 15531 17561
rect 10870 17524 10876 17536
rect 9600 17496 10876 17524
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 11241 17527 11299 17533
rect 11241 17493 11253 17527
rect 11287 17524 11299 17527
rect 12434 17524 12440 17536
rect 11287 17496 12440 17524
rect 11287 17493 11299 17496
rect 11241 17487 11299 17493
rect 12434 17484 12440 17496
rect 12492 17484 12498 17536
rect 14921 17527 14979 17533
rect 14921 17493 14933 17527
rect 14967 17524 14979 17527
rect 15378 17524 15384 17536
rect 14967 17496 15384 17524
rect 14967 17493 14979 17496
rect 14921 17487 14979 17493
rect 15378 17484 15384 17496
rect 15436 17484 15442 17536
rect 1104 17434 17388 17456
rect 1104 17382 3696 17434
rect 3748 17382 3760 17434
rect 3812 17382 3824 17434
rect 3876 17382 3888 17434
rect 3940 17382 9124 17434
rect 9176 17382 9188 17434
rect 9240 17382 9252 17434
rect 9304 17382 9316 17434
rect 9368 17382 14552 17434
rect 14604 17382 14616 17434
rect 14668 17382 14680 17434
rect 14732 17382 14744 17434
rect 14796 17382 17388 17434
rect 1104 17360 17388 17382
rect 3326 17280 3332 17332
rect 3384 17320 3390 17332
rect 6825 17323 6883 17329
rect 3384 17292 6408 17320
rect 3384 17280 3390 17292
rect 5074 17144 5080 17196
rect 5132 17184 5138 17196
rect 5445 17187 5503 17193
rect 5445 17184 5457 17187
rect 5132 17156 5457 17184
rect 5132 17144 5138 17156
rect 5445 17153 5457 17156
rect 5491 17153 5503 17187
rect 5445 17147 5503 17153
rect 2317 17119 2375 17125
rect 2317 17085 2329 17119
rect 2363 17116 2375 17119
rect 2406 17116 2412 17128
rect 2363 17088 2412 17116
rect 2363 17085 2375 17088
rect 2317 17079 2375 17085
rect 2406 17076 2412 17088
rect 2464 17076 2470 17128
rect 4798 17076 4804 17128
rect 4856 17116 4862 17128
rect 5258 17116 5264 17128
rect 4856 17088 4901 17116
rect 5219 17088 5264 17116
rect 4856 17076 4862 17088
rect 5258 17076 5264 17088
rect 5316 17076 5322 17128
rect 5350 17076 5356 17128
rect 5408 17116 5414 17128
rect 5629 17119 5687 17125
rect 5629 17116 5641 17119
rect 5408 17088 5641 17116
rect 5408 17076 5414 17088
rect 5629 17085 5641 17088
rect 5675 17085 5687 17119
rect 6380 17116 6408 17292
rect 6825 17289 6837 17323
rect 6871 17320 6883 17323
rect 7098 17320 7104 17332
rect 6871 17292 7104 17320
rect 6871 17289 6883 17292
rect 6825 17283 6883 17289
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 16393 17323 16451 17329
rect 16393 17320 16405 17323
rect 15620 17292 16405 17320
rect 15620 17280 15626 17292
rect 16393 17289 16405 17292
rect 16439 17289 16451 17323
rect 16393 17283 16451 17289
rect 6730 17212 6736 17264
rect 6788 17252 6794 17264
rect 6788 17224 7972 17252
rect 6788 17212 6794 17224
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17184 7435 17187
rect 7650 17184 7656 17196
rect 7423 17156 7656 17184
rect 7423 17153 7435 17156
rect 7377 17147 7435 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 7944 17193 7972 17224
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17153 7987 17187
rect 7929 17147 7987 17153
rect 10134 17144 10140 17196
rect 10192 17184 10198 17196
rect 10873 17187 10931 17193
rect 10873 17184 10885 17187
rect 10192 17156 10885 17184
rect 10192 17144 10198 17156
rect 10873 17153 10885 17156
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17184 14059 17187
rect 14918 17184 14924 17196
rect 14047 17156 14136 17184
rect 14879 17156 14924 17184
rect 14047 17153 14059 17156
rect 14001 17147 14059 17153
rect 14108 17128 14136 17156
rect 14918 17144 14924 17156
rect 14976 17144 14982 17196
rect 6950 17119 7008 17125
rect 6950 17116 6962 17119
rect 6380 17088 6962 17116
rect 5629 17079 5687 17085
rect 6950 17085 6962 17088
rect 6996 17116 7008 17119
rect 7469 17119 7527 17125
rect 7469 17116 7481 17119
rect 6996 17088 7481 17116
rect 6996 17085 7008 17088
rect 6950 17079 7008 17085
rect 7469 17085 7481 17088
rect 7515 17116 7527 17119
rect 7834 17116 7840 17128
rect 7515 17088 7840 17116
rect 7515 17085 7527 17088
rect 7469 17079 7527 17085
rect 7834 17076 7840 17088
rect 7892 17076 7898 17128
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 10735 17088 12480 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 4430 17048 4436 17060
rect 4094 17020 4436 17048
rect 4430 17008 4436 17020
rect 4488 17008 4494 17060
rect 4522 17008 4528 17060
rect 4580 17048 4586 17060
rect 5534 17048 5540 17060
rect 4580 17020 4625 17048
rect 5495 17020 5540 17048
rect 4580 17008 4586 17020
rect 5534 17008 5540 17020
rect 5592 17008 5598 17060
rect 8202 17048 8208 17060
rect 8163 17020 8208 17048
rect 8202 17008 8208 17020
rect 8260 17008 8266 17060
rect 9490 17048 9496 17060
rect 9430 17020 9496 17048
rect 9490 17008 9496 17020
rect 9548 17008 9554 17060
rect 2501 16983 2559 16989
rect 2501 16949 2513 16983
rect 2547 16980 2559 16983
rect 2866 16980 2872 16992
rect 2547 16952 2872 16980
rect 2547 16949 2559 16952
rect 2501 16943 2559 16949
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 3053 16983 3111 16989
rect 3053 16949 3065 16983
rect 3099 16980 3111 16983
rect 3234 16980 3240 16992
rect 3099 16952 3240 16980
rect 3099 16949 3111 16952
rect 3053 16943 3111 16949
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 5166 16940 5172 16992
rect 5224 16980 5230 16992
rect 5353 16983 5411 16989
rect 5353 16980 5365 16983
rect 5224 16952 5365 16980
rect 5224 16940 5230 16952
rect 5353 16949 5365 16952
rect 5399 16949 5411 16983
rect 5353 16943 5411 16949
rect 7009 16983 7067 16989
rect 7009 16949 7021 16983
rect 7055 16980 7067 16983
rect 7650 16980 7656 16992
rect 7055 16952 7656 16980
rect 7055 16949 7067 16952
rect 7009 16943 7067 16949
rect 7650 16940 7656 16952
rect 7708 16940 7714 16992
rect 7926 16940 7932 16992
rect 7984 16980 7990 16992
rect 9677 16983 9735 16989
rect 9677 16980 9689 16983
rect 7984 16952 9689 16980
rect 7984 16940 7990 16952
rect 9677 16949 9689 16952
rect 9723 16949 9735 16983
rect 10502 16980 10508 16992
rect 10463 16952 10508 16980
rect 9677 16943 9735 16949
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 12250 16980 12256 16992
rect 12211 16952 12256 16980
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 12452 16980 12480 17088
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 14645 17119 14703 17125
rect 14645 17116 14657 17119
rect 14148 17088 14657 17116
rect 14148 17076 14154 17088
rect 14645 17085 14657 17088
rect 14691 17085 14703 17119
rect 14645 17079 14703 17085
rect 13170 17008 13176 17060
rect 13228 17008 13234 17060
rect 13722 17048 13728 17060
rect 13683 17020 13728 17048
rect 13722 17008 13728 17020
rect 13780 17008 13786 17060
rect 15930 17008 15936 17060
rect 15988 17008 15994 17060
rect 15286 16980 15292 16992
rect 12452 16952 15292 16980
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 1104 16890 17388 16912
rect 1104 16838 6410 16890
rect 6462 16838 6474 16890
rect 6526 16838 6538 16890
rect 6590 16838 6602 16890
rect 6654 16838 11838 16890
rect 11890 16838 11902 16890
rect 11954 16838 11966 16890
rect 12018 16838 12030 16890
rect 12082 16838 17388 16890
rect 1104 16816 17388 16838
rect 2777 16779 2835 16785
rect 2777 16745 2789 16779
rect 2823 16776 2835 16779
rect 3326 16776 3332 16788
rect 2823 16748 3332 16776
rect 2823 16745 2835 16748
rect 2777 16739 2835 16745
rect 3326 16736 3332 16748
rect 3384 16736 3390 16788
rect 6641 16779 6699 16785
rect 6641 16745 6653 16779
rect 6687 16776 6699 16779
rect 7190 16776 7196 16788
rect 6687 16748 7196 16776
rect 6687 16745 6699 16748
rect 6641 16739 6699 16745
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 8202 16776 8208 16788
rect 8163 16748 8208 16776
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 9766 16736 9772 16788
rect 9824 16776 9830 16788
rect 9953 16779 10011 16785
rect 9953 16776 9965 16779
rect 9824 16748 9965 16776
rect 9824 16736 9830 16748
rect 9953 16745 9965 16748
rect 9999 16745 10011 16779
rect 9953 16739 10011 16745
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16776 10195 16779
rect 10410 16776 10416 16788
rect 10183 16748 10416 16776
rect 10183 16745 10195 16748
rect 10137 16739 10195 16745
rect 10410 16736 10416 16748
rect 10468 16736 10474 16788
rect 12069 16779 12127 16785
rect 12069 16745 12081 16779
rect 12115 16776 12127 16779
rect 12434 16776 12440 16788
rect 12115 16748 12440 16776
rect 12115 16745 12127 16748
rect 12069 16739 12127 16745
rect 12434 16736 12440 16748
rect 12492 16736 12498 16788
rect 13170 16776 13176 16788
rect 13131 16748 13176 16776
rect 13170 16736 13176 16748
rect 13228 16736 13234 16788
rect 13630 16776 13636 16788
rect 13591 16748 13636 16776
rect 13630 16736 13636 16748
rect 13688 16736 13694 16788
rect 15197 16779 15255 16785
rect 15197 16776 15209 16779
rect 14844 16748 15209 16776
rect 5166 16708 5172 16720
rect 5127 16680 5172 16708
rect 5166 16668 5172 16680
rect 5224 16668 5230 16720
rect 5902 16668 5908 16720
rect 5960 16668 5966 16720
rect 7926 16708 7932 16720
rect 7887 16680 7932 16708
rect 7926 16668 7932 16680
rect 7984 16668 7990 16720
rect 13354 16708 13360 16720
rect 11256 16680 13360 16708
rect 2774 16643 2832 16649
rect 2774 16609 2786 16643
rect 2820 16640 2832 16643
rect 2820 16612 3280 16640
rect 2820 16609 2832 16612
rect 2774 16603 2832 16609
rect 3252 16584 3280 16612
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 4798 16640 4804 16652
rect 4212 16612 4804 16640
rect 4212 16600 4218 16612
rect 4798 16600 4804 16612
rect 4856 16640 4862 16652
rect 4893 16643 4951 16649
rect 4893 16640 4905 16643
rect 4856 16612 4905 16640
rect 4856 16600 4862 16612
rect 4893 16609 4905 16612
rect 4939 16609 4951 16643
rect 7650 16640 7656 16652
rect 7611 16612 7656 16640
rect 4893 16603 4951 16609
rect 7650 16600 7656 16612
rect 7708 16600 7714 16652
rect 7834 16640 7840 16652
rect 7795 16612 7840 16640
rect 7834 16600 7840 16612
rect 7892 16600 7898 16652
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16640 8079 16643
rect 8202 16640 8208 16652
rect 8067 16612 8208 16640
rect 8067 16609 8079 16612
rect 8021 16603 8079 16609
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 9950 16600 9956 16652
rect 10008 16640 10014 16652
rect 10078 16643 10136 16649
rect 10078 16640 10090 16643
rect 10008 16612 10090 16640
rect 10008 16600 10014 16612
rect 10078 16609 10090 16612
rect 10124 16640 10136 16643
rect 10502 16640 10508 16652
rect 10124 16612 10508 16640
rect 10124 16609 10136 16612
rect 10078 16603 10136 16609
rect 10502 16600 10508 16612
rect 10560 16640 10566 16652
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 10560 16612 10609 16640
rect 10560 16600 10566 16612
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 11256 16649 11284 16680
rect 13354 16668 13360 16680
rect 13412 16668 13418 16720
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 10744 16612 11161 16640
rect 10744 16600 10750 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 12066 16643 12124 16649
rect 12066 16609 12078 16643
rect 12112 16640 12124 16643
rect 12250 16640 12256 16652
rect 12112 16612 12256 16640
rect 12112 16609 12124 16612
rect 12066 16603 12124 16609
rect 12250 16600 12256 16612
rect 12308 16640 12314 16652
rect 12529 16643 12587 16649
rect 12529 16640 12541 16643
rect 12308 16612 12541 16640
rect 12308 16600 12314 16612
rect 12529 16609 12541 16612
rect 12575 16609 12587 16643
rect 12529 16603 12587 16609
rect 12989 16643 13047 16649
rect 12989 16609 13001 16643
rect 13035 16640 13047 16643
rect 13262 16640 13268 16652
rect 13035 16612 13268 16640
rect 13035 16609 13047 16612
rect 12989 16603 13047 16609
rect 13262 16600 13268 16612
rect 13320 16640 13326 16652
rect 14844 16649 14872 16748
rect 15197 16745 15209 16748
rect 15243 16776 15255 16779
rect 15378 16776 15384 16788
rect 15243 16748 15384 16776
rect 15243 16745 15255 16748
rect 15197 16739 15255 16745
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 15930 16776 15936 16788
rect 15891 16748 15936 16776
rect 15930 16736 15936 16748
rect 15988 16736 15994 16788
rect 13817 16643 13875 16649
rect 13817 16640 13829 16643
rect 13320 16612 13829 16640
rect 13320 16600 13326 16612
rect 13817 16609 13829 16612
rect 13863 16640 13875 16643
rect 14737 16643 14795 16649
rect 13863 16612 14688 16640
rect 13863 16609 13875 16612
rect 13817 16603 13875 16609
rect 3234 16572 3240 16584
rect 3195 16544 3240 16572
rect 3234 16532 3240 16544
rect 3292 16532 3298 16584
rect 12434 16572 12440 16584
rect 12395 16544 12440 16572
rect 12434 16532 12440 16544
rect 12492 16532 12498 16584
rect 1486 16464 1492 16516
rect 1544 16504 1550 16516
rect 11885 16507 11943 16513
rect 1544 16476 5028 16504
rect 1544 16464 1550 16476
rect 2590 16436 2596 16448
rect 2551 16408 2596 16436
rect 2590 16396 2596 16408
rect 2648 16396 2654 16448
rect 3145 16439 3203 16445
rect 3145 16405 3157 16439
rect 3191 16436 3203 16439
rect 3326 16436 3332 16448
rect 3191 16408 3332 16436
rect 3191 16405 3203 16408
rect 3145 16399 3203 16405
rect 3326 16396 3332 16408
rect 3384 16396 3390 16448
rect 5000 16436 5028 16476
rect 11885 16473 11897 16507
rect 11931 16504 11943 16507
rect 12066 16504 12072 16516
rect 11931 16476 12072 16504
rect 11931 16473 11943 16476
rect 11885 16467 11943 16473
rect 12066 16464 12072 16476
rect 12124 16504 12130 16516
rect 12342 16504 12348 16516
rect 12124 16476 12348 16504
rect 12124 16464 12130 16476
rect 12342 16464 12348 16476
rect 12400 16464 12406 16516
rect 14660 16504 14688 16612
rect 14737 16609 14749 16643
rect 14783 16609 14795 16643
rect 14737 16603 14795 16609
rect 14829 16643 14887 16649
rect 14829 16609 14841 16643
rect 14875 16609 14887 16643
rect 15194 16640 15200 16652
rect 14829 16603 14887 16609
rect 14936 16612 15200 16640
rect 14752 16572 14780 16603
rect 14936 16572 14964 16612
rect 15194 16600 15200 16612
rect 15252 16640 15258 16652
rect 16114 16640 16120 16652
rect 15252 16612 15297 16640
rect 16075 16612 16120 16640
rect 15252 16600 15258 16612
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 14752 16544 14964 16572
rect 16114 16504 16120 16516
rect 14660 16476 16120 16504
rect 16114 16464 16120 16476
rect 16172 16464 16178 16516
rect 10134 16436 10140 16448
rect 5000 16408 10140 16436
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 10410 16396 10416 16448
rect 10468 16436 10474 16448
rect 10505 16439 10563 16445
rect 10505 16436 10517 16439
rect 10468 16408 10517 16436
rect 10468 16396 10474 16408
rect 10505 16405 10517 16408
rect 10551 16405 10563 16439
rect 10505 16399 10563 16405
rect 15194 16396 15200 16448
rect 15252 16436 15258 16448
rect 15381 16439 15439 16445
rect 15381 16436 15393 16439
rect 15252 16408 15393 16436
rect 15252 16396 15258 16408
rect 15381 16405 15393 16408
rect 15427 16405 15439 16439
rect 15381 16399 15439 16405
rect 1104 16346 17388 16368
rect 1104 16294 3696 16346
rect 3748 16294 3760 16346
rect 3812 16294 3824 16346
rect 3876 16294 3888 16346
rect 3940 16294 9124 16346
rect 9176 16294 9188 16346
rect 9240 16294 9252 16346
rect 9304 16294 9316 16346
rect 9368 16294 14552 16346
rect 14604 16294 14616 16346
rect 14668 16294 14680 16346
rect 14732 16294 14744 16346
rect 14796 16294 17388 16346
rect 1104 16272 17388 16294
rect 2409 16235 2467 16241
rect 2409 16201 2421 16235
rect 2455 16232 2467 16235
rect 2590 16232 2596 16244
rect 2455 16204 2596 16232
rect 2455 16201 2467 16204
rect 2409 16195 2467 16201
rect 2590 16192 2596 16204
rect 2648 16232 2654 16244
rect 4430 16232 4436 16244
rect 2648 16204 4016 16232
rect 4391 16204 4436 16232
rect 2648 16192 2654 16204
rect 2961 16167 3019 16173
rect 2961 16133 2973 16167
rect 3007 16164 3019 16167
rect 3007 16136 3924 16164
rect 3007 16133 3019 16136
rect 2961 16127 3019 16133
rect 1486 16096 1492 16108
rect 1447 16068 1492 16096
rect 1486 16056 1492 16068
rect 1544 16056 1550 16108
rect 2317 16099 2375 16105
rect 2317 16065 2329 16099
rect 2363 16096 2375 16099
rect 2498 16096 2504 16108
rect 2363 16068 2504 16096
rect 2363 16065 2375 16068
rect 2317 16059 2375 16065
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 3160 16068 3832 16096
rect 1670 16028 1676 16040
rect 1631 16000 1676 16028
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 2516 16028 2544 16056
rect 2836 16031 2894 16037
rect 2836 16028 2848 16031
rect 2516 16000 2848 16028
rect 2836 15997 2848 16000
rect 2882 16028 2894 16031
rect 3160 16028 3188 16068
rect 2882 16000 3188 16028
rect 2882 15997 2894 16000
rect 2836 15991 2894 15997
rect 3326 15988 3332 16040
rect 3384 16028 3390 16040
rect 3804 16037 3832 16068
rect 3605 16031 3663 16037
rect 3605 16028 3617 16031
rect 3384 16000 3617 16028
rect 3384 15988 3390 16000
rect 3605 15997 3617 16000
rect 3651 15997 3663 16031
rect 3605 15991 3663 15997
rect 3789 16031 3847 16037
rect 3789 15997 3801 16031
rect 3835 15997 3847 16031
rect 3789 15991 3847 15997
rect 3234 15920 3240 15972
rect 3292 15960 3298 15972
rect 3697 15963 3755 15969
rect 3697 15960 3709 15963
rect 3292 15932 3709 15960
rect 3292 15920 3298 15932
rect 3697 15929 3709 15932
rect 3743 15929 3755 15963
rect 3896 15960 3924 16136
rect 3988 16037 4016 16204
rect 4430 16192 4436 16204
rect 4488 16192 4494 16244
rect 5902 16232 5908 16244
rect 5863 16204 5908 16232
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 7650 16232 7656 16244
rect 7611 16204 7656 16232
rect 7650 16192 7656 16204
rect 7708 16192 7714 16244
rect 8754 16232 8760 16244
rect 8715 16204 8760 16232
rect 8754 16192 8760 16204
rect 8812 16192 8818 16244
rect 9401 16235 9459 16241
rect 9401 16201 9413 16235
rect 9447 16232 9459 16235
rect 9490 16232 9496 16244
rect 9447 16204 9496 16232
rect 9447 16201 9459 16204
rect 9401 16195 9459 16201
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 12621 16235 12679 16241
rect 12621 16201 12633 16235
rect 12667 16232 12679 16235
rect 13722 16232 13728 16244
rect 12667 16204 13728 16232
rect 12667 16201 12679 16204
rect 12621 16195 12679 16201
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 15286 16232 15292 16244
rect 15247 16204 15292 16232
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 7193 16167 7251 16173
rect 7193 16133 7205 16167
rect 7239 16164 7251 16167
rect 9858 16164 9864 16176
rect 7239 16136 9864 16164
rect 7239 16133 7251 16136
rect 7193 16127 7251 16133
rect 9858 16124 9864 16136
rect 9916 16124 9922 16176
rect 7926 16056 7932 16108
rect 7984 16096 7990 16108
rect 8297 16099 8355 16105
rect 8297 16096 8309 16099
rect 7984 16068 8309 16096
rect 7984 16056 7990 16068
rect 8297 16065 8309 16068
rect 8343 16065 8355 16099
rect 16574 16096 16580 16108
rect 8297 16059 8355 16065
rect 10888 16068 11100 16096
rect 3973 16031 4031 16037
rect 3973 15997 3985 16031
rect 4019 15997 4031 16031
rect 4614 16028 4620 16040
rect 4527 16000 4620 16028
rect 3973 15991 4031 15997
rect 4614 15988 4620 16000
rect 4672 16028 4678 16040
rect 5721 16031 5779 16037
rect 5721 16028 5733 16031
rect 4672 16000 5733 16028
rect 4672 15988 4678 16000
rect 5721 15997 5733 16000
rect 5767 15997 5779 16031
rect 5721 15991 5779 15997
rect 7009 16031 7067 16037
rect 7009 15997 7021 16031
rect 7055 15997 7067 16031
rect 7009 15991 7067 15997
rect 7834 16031 7892 16037
rect 7834 15997 7846 16031
rect 7880 16028 7892 16031
rect 7944 16028 7972 16056
rect 8202 16028 8208 16040
rect 7880 16000 7972 16028
rect 8163 16000 8208 16028
rect 7880 15997 7892 16000
rect 7834 15991 7892 15997
rect 4430 15960 4436 15972
rect 3896 15932 4436 15960
rect 3697 15923 3755 15929
rect 4430 15920 4436 15932
rect 4488 15920 4494 15972
rect 1857 15895 1915 15901
rect 1857 15861 1869 15895
rect 1903 15892 1915 15895
rect 2038 15892 2044 15904
rect 1903 15864 2044 15892
rect 1903 15861 1915 15864
rect 1857 15855 1915 15861
rect 2038 15852 2044 15864
rect 2096 15852 2102 15904
rect 2590 15852 2596 15904
rect 2648 15892 2654 15904
rect 2777 15895 2835 15901
rect 2777 15892 2789 15895
rect 2648 15864 2789 15892
rect 2648 15852 2654 15864
rect 2777 15861 2789 15864
rect 2823 15861 2835 15895
rect 2777 15855 2835 15861
rect 3421 15895 3479 15901
rect 3421 15861 3433 15895
rect 3467 15892 3479 15895
rect 4522 15892 4528 15904
rect 3467 15864 4528 15892
rect 3467 15861 3479 15864
rect 3421 15855 3479 15861
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 5736 15892 5764 15991
rect 7024 15960 7052 15991
rect 8202 15988 8208 16000
rect 8260 15988 8266 16040
rect 8938 16028 8944 16040
rect 8899 16000 8944 16028
rect 8938 15988 8944 16000
rect 8996 16028 9002 16040
rect 9585 16031 9643 16037
rect 9585 16028 9597 16031
rect 8996 16000 9597 16028
rect 8996 15988 9002 16000
rect 9585 15997 9597 16000
rect 9631 15997 9643 16031
rect 9585 15991 9643 15997
rect 10594 16031 10652 16037
rect 10594 15997 10606 16031
rect 10640 16028 10652 16031
rect 10888 16028 10916 16068
rect 11072 16037 11100 16068
rect 15488 16068 16580 16096
rect 10640 16000 10916 16028
rect 10965 16031 11023 16037
rect 10640 15997 10652 16000
rect 10594 15991 10652 15997
rect 10965 15997 10977 16031
rect 11011 15997 11023 16031
rect 10965 15991 11023 15997
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 16028 11115 16031
rect 11238 16028 11244 16040
rect 11103 16000 11244 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 9674 15960 9680 15972
rect 7024 15932 9680 15960
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 7098 15892 7104 15904
rect 5736 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 7837 15895 7895 15901
rect 7837 15861 7849 15895
rect 7883 15892 7895 15895
rect 8202 15892 8208 15904
rect 7883 15864 8208 15892
rect 7883 15861 7895 15864
rect 7837 15855 7895 15861
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10410 15892 10416 15904
rect 9916 15864 10416 15892
rect 9916 15852 9922 15864
rect 10410 15852 10416 15864
rect 10468 15852 10474 15904
rect 10594 15892 10600 15904
rect 10507 15864 10600 15892
rect 10594 15852 10600 15864
rect 10652 15892 10658 15904
rect 10980 15892 11008 15991
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 12066 16028 12072 16040
rect 12027 16000 12072 16028
rect 12066 15988 12072 16000
rect 12124 15988 12130 16040
rect 12158 15988 12164 16040
rect 12216 16028 12222 16040
rect 12253 16031 12311 16037
rect 12253 16028 12265 16031
rect 12216 16000 12265 16028
rect 12216 15988 12222 16000
rect 12253 15997 12265 16000
rect 12299 15997 12311 16031
rect 12434 16028 12440 16040
rect 12395 16000 12440 16028
rect 12253 15991 12311 15997
rect 12434 15988 12440 16000
rect 12492 15988 12498 16040
rect 13262 16028 13268 16040
rect 13223 16000 13268 16028
rect 13262 15988 13268 16000
rect 13320 15988 13326 16040
rect 13906 16028 13912 16040
rect 13867 16000 13912 16028
rect 13906 15988 13912 16000
rect 13964 15988 13970 16040
rect 14277 16031 14335 16037
rect 14277 15997 14289 16031
rect 14323 16028 14335 16031
rect 15010 16028 15016 16040
rect 14323 16000 15016 16028
rect 14323 15997 14335 16000
rect 14277 15991 14335 15997
rect 15010 15988 15016 16000
rect 15068 15988 15074 16040
rect 15488 16037 15516 16068
rect 16574 16056 16580 16068
rect 16632 16056 16638 16108
rect 15473 16031 15531 16037
rect 15473 15997 15485 16031
rect 15519 15997 15531 16031
rect 15473 15991 15531 15997
rect 15933 16031 15991 16037
rect 15933 15997 15945 16031
rect 15979 16028 15991 16031
rect 16114 16028 16120 16040
rect 15979 16000 16120 16028
rect 15979 15997 15991 16000
rect 15933 15991 15991 15997
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 12342 15960 12348 15972
rect 12303 15932 12348 15960
rect 12342 15920 12348 15932
rect 12400 15920 12406 15972
rect 14090 15960 14096 15972
rect 14051 15932 14096 15960
rect 14090 15920 14096 15932
rect 14148 15920 14154 15972
rect 14185 15963 14243 15969
rect 14185 15929 14197 15963
rect 14231 15960 14243 15963
rect 14918 15960 14924 15972
rect 14231 15932 14924 15960
rect 14231 15929 14243 15932
rect 14185 15923 14243 15929
rect 14918 15920 14924 15932
rect 14976 15920 14982 15972
rect 10652 15864 11008 15892
rect 10652 15852 10658 15864
rect 12710 15852 12716 15904
rect 12768 15892 12774 15904
rect 13081 15895 13139 15901
rect 13081 15892 13093 15895
rect 12768 15864 13093 15892
rect 12768 15852 12774 15864
rect 13081 15861 13093 15864
rect 13127 15861 13139 15895
rect 13081 15855 13139 15861
rect 14274 15852 14280 15904
rect 14332 15892 14338 15904
rect 14461 15895 14519 15901
rect 14461 15892 14473 15895
rect 14332 15864 14473 15892
rect 14332 15852 14338 15864
rect 14461 15861 14473 15864
rect 14507 15861 14519 15895
rect 14461 15855 14519 15861
rect 16117 15895 16175 15901
rect 16117 15861 16129 15895
rect 16163 15892 16175 15895
rect 16206 15892 16212 15904
rect 16163 15864 16212 15892
rect 16163 15861 16175 15864
rect 16117 15855 16175 15861
rect 16206 15852 16212 15864
rect 16264 15852 16270 15904
rect 1104 15802 17388 15824
rect 1104 15750 6410 15802
rect 6462 15750 6474 15802
rect 6526 15750 6538 15802
rect 6590 15750 6602 15802
rect 6654 15750 11838 15802
rect 11890 15750 11902 15802
rect 11954 15750 11966 15802
rect 12018 15750 12030 15802
rect 12082 15750 17388 15802
rect 1104 15728 17388 15750
rect 2041 15691 2099 15697
rect 2041 15657 2053 15691
rect 2087 15688 2099 15691
rect 2087 15660 2452 15688
rect 2087 15657 2099 15660
rect 2041 15651 2099 15657
rect 2424 15561 2452 15660
rect 5534 15648 5540 15700
rect 5592 15688 5598 15700
rect 5997 15691 6055 15697
rect 5997 15688 6009 15691
rect 5592 15660 6009 15688
rect 5592 15648 5598 15660
rect 5997 15657 6009 15660
rect 6043 15657 6055 15691
rect 5997 15651 6055 15657
rect 10413 15691 10471 15697
rect 10413 15657 10425 15691
rect 10459 15688 10471 15691
rect 10459 15660 11192 15688
rect 10459 15657 10471 15660
rect 10413 15651 10471 15657
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 11164 15629 11192 15660
rect 11238 15648 11244 15700
rect 11296 15688 11302 15700
rect 12621 15691 12679 15697
rect 12621 15688 12633 15691
rect 11296 15660 12633 15688
rect 11296 15648 11302 15660
rect 12621 15657 12633 15660
rect 12667 15657 12679 15691
rect 13262 15688 13268 15700
rect 13223 15660 13268 15688
rect 12621 15651 12679 15657
rect 13262 15648 13268 15660
rect 13320 15648 13326 15700
rect 10045 15623 10103 15629
rect 10045 15620 10057 15623
rect 10008 15592 10057 15620
rect 10008 15580 10014 15592
rect 10045 15589 10057 15592
rect 10091 15589 10103 15623
rect 10045 15583 10103 15589
rect 11149 15623 11207 15629
rect 11149 15589 11161 15623
rect 11195 15589 11207 15623
rect 12710 15620 12716 15632
rect 12374 15592 12716 15620
rect 11149 15583 11207 15589
rect 12710 15580 12716 15592
rect 12768 15580 12774 15632
rect 15194 15620 15200 15632
rect 15155 15592 15200 15620
rect 15194 15580 15200 15592
rect 15252 15580 15258 15632
rect 16206 15580 16212 15632
rect 16264 15580 16270 15632
rect 2038 15555 2096 15561
rect 2038 15521 2050 15555
rect 2084 15552 2096 15555
rect 2409 15555 2467 15561
rect 2084 15524 2268 15552
rect 2084 15521 2096 15524
rect 2038 15515 2096 15521
rect 2240 15496 2268 15524
rect 2409 15521 2421 15555
rect 2455 15552 2467 15555
rect 2958 15552 2964 15564
rect 2455 15524 2964 15552
rect 2455 15521 2467 15524
rect 2409 15515 2467 15521
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 4614 15552 4620 15564
rect 4479 15524 4620 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 5994 15512 6000 15564
rect 6052 15552 6058 15564
rect 6181 15555 6239 15561
rect 6181 15552 6193 15555
rect 6052 15524 6193 15552
rect 6052 15512 6058 15524
rect 6181 15521 6193 15524
rect 6227 15521 6239 15555
rect 6181 15515 6239 15521
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15552 6699 15555
rect 6822 15552 6828 15564
rect 6687 15524 6828 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 6822 15512 6828 15524
rect 6880 15512 6886 15564
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 7285 15555 7343 15561
rect 7285 15552 7297 15555
rect 7156 15524 7297 15552
rect 7156 15512 7162 15524
rect 7285 15521 7297 15524
rect 7331 15521 7343 15555
rect 8110 15552 8116 15564
rect 8071 15524 8116 15552
rect 7285 15515 7343 15521
rect 2222 15444 2228 15496
rect 2280 15484 2286 15496
rect 2501 15487 2559 15493
rect 2501 15484 2513 15487
rect 2280 15456 2513 15484
rect 2280 15444 2286 15456
rect 2501 15453 2513 15456
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 7300 15416 7328 15515
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 9858 15552 9864 15564
rect 9819 15524 9864 15552
rect 9858 15512 9864 15524
rect 9916 15512 9922 15564
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15521 10195 15555
rect 10137 15515 10195 15521
rect 10229 15555 10287 15561
rect 10229 15521 10241 15555
rect 10275 15552 10287 15555
rect 10594 15552 10600 15564
rect 10275 15524 10600 15552
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 10152 15484 10180 15515
rect 10594 15512 10600 15524
rect 10652 15512 10658 15564
rect 10870 15552 10876 15564
rect 10831 15524 10876 15552
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15552 13139 15555
rect 13354 15552 13360 15564
rect 13127 15524 13360 15552
rect 13127 15521 13139 15524
rect 13081 15515 13139 15521
rect 13354 15512 13360 15524
rect 13412 15512 13418 15564
rect 11238 15484 11244 15496
rect 10152 15456 11244 15484
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 13998 15444 14004 15496
rect 14056 15484 14062 15496
rect 14921 15487 14979 15493
rect 14921 15484 14933 15487
rect 14056 15456 14933 15484
rect 14056 15444 14062 15456
rect 14921 15453 14933 15456
rect 14967 15453 14979 15487
rect 14921 15447 14979 15453
rect 7929 15419 7987 15425
rect 7929 15416 7941 15419
rect 7300 15388 7941 15416
rect 7929 15385 7941 15388
rect 7975 15385 7987 15419
rect 7929 15379 7987 15385
rect 1854 15348 1860 15360
rect 1815 15320 1860 15348
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 4614 15348 4620 15360
rect 4575 15320 4620 15348
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 6730 15308 6736 15360
rect 6788 15348 6794 15360
rect 6825 15351 6883 15357
rect 6825 15348 6837 15351
rect 6788 15320 6837 15348
rect 6788 15308 6794 15320
rect 6825 15317 6837 15320
rect 6871 15317 6883 15351
rect 6825 15311 6883 15317
rect 7469 15351 7527 15357
rect 7469 15317 7481 15351
rect 7515 15348 7527 15351
rect 7558 15348 7564 15360
rect 7515 15320 7564 15348
rect 7515 15317 7527 15320
rect 7469 15311 7527 15317
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 15010 15308 15016 15360
rect 15068 15348 15074 15360
rect 16669 15351 16727 15357
rect 16669 15348 16681 15351
rect 15068 15320 16681 15348
rect 15068 15308 15074 15320
rect 16669 15317 16681 15320
rect 16715 15317 16727 15351
rect 16669 15311 16727 15317
rect 1104 15258 17388 15280
rect 1104 15206 3696 15258
rect 3748 15206 3760 15258
rect 3812 15206 3824 15258
rect 3876 15206 3888 15258
rect 3940 15206 9124 15258
rect 9176 15206 9188 15258
rect 9240 15206 9252 15258
rect 9304 15206 9316 15258
rect 9368 15206 14552 15258
rect 14604 15206 14616 15258
rect 14668 15206 14680 15258
rect 14732 15206 14744 15258
rect 14796 15206 17388 15258
rect 1104 15184 17388 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1765 15147 1823 15153
rect 1765 15144 1777 15147
rect 1728 15116 1777 15144
rect 1728 15104 1734 15116
rect 1765 15113 1777 15116
rect 1811 15113 1823 15147
rect 1765 15107 1823 15113
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 6730 15144 6736 15156
rect 4212 15116 6736 15144
rect 4212 15104 4218 15116
rect 6730 15104 6736 15116
rect 6788 15144 6794 15156
rect 6788 15116 6868 15144
rect 6788 15104 6794 15116
rect 5261 15079 5319 15085
rect 5261 15045 5273 15079
rect 5307 15076 5319 15079
rect 5534 15076 5540 15088
rect 5307 15048 5540 15076
rect 5307 15045 5319 15048
rect 5261 15039 5319 15045
rect 5534 15036 5540 15048
rect 5592 15036 5598 15088
rect 6840 15017 6868 15116
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 8573 15147 8631 15153
rect 8573 15144 8585 15147
rect 8260 15116 8585 15144
rect 8260 15104 8266 15116
rect 8573 15113 8585 15116
rect 8619 15113 8631 15147
rect 8573 15107 8631 15113
rect 10594 15104 10600 15156
rect 10652 15144 10658 15156
rect 10781 15147 10839 15153
rect 10781 15144 10793 15147
rect 10652 15116 10793 15144
rect 10652 15104 10658 15116
rect 10781 15113 10793 15116
rect 10827 15113 10839 15147
rect 10781 15107 10839 15113
rect 10870 15104 10876 15156
rect 10928 15144 10934 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 10928 15116 11529 15144
rect 10928 15104 10934 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 13265 15147 13323 15153
rect 13265 15113 13277 15147
rect 13311 15144 13323 15147
rect 14090 15144 14096 15156
rect 13311 15116 14096 15144
rect 13311 15113 13323 15116
rect 13265 15107 13323 15113
rect 6825 15011 6883 15017
rect 5644 14980 5948 15008
rect 1946 14940 1952 14952
rect 1907 14912 1952 14940
rect 1946 14900 1952 14912
rect 2004 14900 2010 14952
rect 3970 14900 3976 14952
rect 4028 14940 4034 14952
rect 4028 14912 4073 14940
rect 4028 14900 4034 14912
rect 4338 14900 4344 14952
rect 4396 14940 4402 14952
rect 4617 14943 4675 14949
rect 4617 14940 4629 14943
rect 4396 14912 4629 14940
rect 4396 14900 4402 14912
rect 4617 14909 4629 14912
rect 4663 14909 4675 14943
rect 4617 14903 4675 14909
rect 5442 14943 5500 14949
rect 5442 14909 5454 14943
rect 5488 14940 5500 14943
rect 5644 14940 5672 14980
rect 5810 14940 5816 14952
rect 5488 14912 5672 14940
rect 5771 14912 5816 14940
rect 5488 14909 5500 14912
rect 5442 14903 5500 14909
rect 5810 14900 5816 14912
rect 5868 14900 5874 14952
rect 5920 14949 5948 14980
rect 6825 14977 6837 15011
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 9033 15011 9091 15017
rect 9033 14977 9045 15011
rect 9079 15008 9091 15011
rect 9674 15008 9680 15020
rect 9079 14980 9680 15008
rect 9079 14977 9091 14980
rect 9033 14971 9091 14977
rect 9674 14968 9680 14980
rect 9732 15008 9738 15020
rect 10870 15008 10876 15020
rect 9732 14980 10876 15008
rect 9732 14968 9738 14980
rect 10870 14968 10876 14980
rect 10928 14968 10934 15020
rect 5905 14943 5963 14949
rect 5905 14909 5917 14943
rect 5951 14940 5963 14943
rect 6730 14940 6736 14952
rect 5951 14912 6736 14940
rect 5951 14909 5963 14912
rect 5905 14903 5963 14909
rect 6730 14900 6736 14912
rect 6788 14900 6794 14952
rect 11330 14940 11336 14952
rect 11291 14912 11336 14940
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 3694 14872 3700 14884
rect 2222 14804 2228 14816
rect 2183 14776 2228 14804
rect 2222 14764 2228 14776
rect 2280 14764 2286 14816
rect 3252 14804 3280 14858
rect 3655 14844 3700 14872
rect 3694 14832 3700 14844
rect 3752 14832 3758 14884
rect 5718 14832 5724 14884
rect 5776 14872 5782 14884
rect 7101 14875 7159 14881
rect 7101 14872 7113 14875
rect 5776 14844 7113 14872
rect 5776 14832 5782 14844
rect 7101 14841 7113 14844
rect 7147 14841 7159 14875
rect 7101 14835 7159 14841
rect 7558 14832 7564 14884
rect 7616 14832 7622 14884
rect 9309 14875 9367 14881
rect 9309 14841 9321 14875
rect 9355 14841 9367 14875
rect 9309 14835 9367 14841
rect 4433 14807 4491 14813
rect 4433 14804 4445 14807
rect 3252 14776 4445 14804
rect 4433 14773 4445 14776
rect 4479 14773 4491 14807
rect 4433 14767 4491 14773
rect 5445 14807 5503 14813
rect 5445 14773 5457 14807
rect 5491 14804 5503 14807
rect 5810 14804 5816 14816
rect 5491 14776 5816 14804
rect 5491 14773 5503 14776
rect 5445 14767 5503 14773
rect 5810 14764 5816 14776
rect 5868 14764 5874 14816
rect 5994 14764 6000 14816
rect 6052 14804 6058 14816
rect 9324 14804 9352 14835
rect 9766 14832 9772 14884
rect 9824 14832 9830 14884
rect 11532 14872 11560 15107
rect 14090 15104 14096 15116
rect 14148 15104 14154 15156
rect 13814 15076 13820 15088
rect 12406 15048 13820 15076
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12406 14940 12434 15048
rect 13814 15036 13820 15048
rect 13872 15036 13878 15088
rect 14093 15011 14151 15017
rect 13004 14980 13860 15008
rect 12299 14912 12434 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12802 14900 12808 14952
rect 12860 14940 12866 14952
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12860 14912 12909 14940
rect 12860 14900 12866 14912
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 13004 14884 13032 14980
rect 13832 14952 13860 14980
rect 14093 14977 14105 15011
rect 14139 15008 14151 15011
rect 14182 15008 14188 15020
rect 14139 14980 14188 15008
rect 14139 14977 14151 14980
rect 14093 14971 14151 14977
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 14826 14968 14832 15020
rect 14884 15008 14890 15020
rect 15470 15008 15476 15020
rect 14884 14980 15476 15008
rect 14884 14968 14890 14980
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14909 13139 14943
rect 13814 14940 13820 14952
rect 13727 14912 13820 14940
rect 13081 14903 13139 14909
rect 12986 14872 12992 14884
rect 11532 14844 12992 14872
rect 12986 14832 12992 14844
rect 13044 14832 13050 14884
rect 13096 14872 13124 14903
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 16390 14940 16396 14952
rect 16351 14912 16396 14940
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 13096 14844 14320 14872
rect 6052 14776 9352 14804
rect 12437 14807 12495 14813
rect 6052 14764 6058 14776
rect 12437 14773 12449 14807
rect 12483 14804 12495 14807
rect 13170 14804 13176 14816
rect 12483 14776 13176 14804
rect 12483 14773 12495 14776
rect 12437 14767 12495 14773
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 13998 14804 14004 14816
rect 13872 14776 14004 14804
rect 13872 14764 13878 14776
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 14292 14804 14320 14844
rect 14366 14832 14372 14884
rect 14424 14872 14430 14884
rect 14424 14844 14582 14872
rect 14424 14832 14430 14844
rect 14826 14804 14832 14816
rect 14292 14776 14832 14804
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 14918 14764 14924 14816
rect 14976 14804 14982 14816
rect 15565 14807 15623 14813
rect 15565 14804 15577 14807
rect 14976 14776 15577 14804
rect 14976 14764 14982 14776
rect 15565 14773 15577 14776
rect 15611 14773 15623 14807
rect 15565 14767 15623 14773
rect 16114 14764 16120 14816
rect 16172 14804 16178 14816
rect 16209 14807 16267 14813
rect 16209 14804 16221 14807
rect 16172 14776 16221 14804
rect 16172 14764 16178 14776
rect 16209 14773 16221 14776
rect 16255 14773 16267 14807
rect 16209 14767 16267 14773
rect 1104 14714 17388 14736
rect 1104 14662 6410 14714
rect 6462 14662 6474 14714
rect 6526 14662 6538 14714
rect 6590 14662 6602 14714
rect 6654 14662 11838 14714
rect 11890 14662 11902 14714
rect 11954 14662 11966 14714
rect 12018 14662 12030 14714
rect 12082 14662 17388 14714
rect 1104 14640 17388 14662
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 1949 14603 2007 14609
rect 1949 14600 1961 14603
rect 1912 14572 1961 14600
rect 1912 14560 1918 14572
rect 1949 14569 1961 14572
rect 1995 14569 2007 14603
rect 1949 14563 2007 14569
rect 3145 14603 3203 14609
rect 3145 14569 3157 14603
rect 3191 14600 3203 14603
rect 3694 14600 3700 14612
rect 3191 14572 3700 14600
rect 3191 14569 3203 14572
rect 3145 14563 3203 14569
rect 3694 14560 3700 14572
rect 3752 14560 3758 14612
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 5868 14572 6009 14600
rect 5868 14560 5874 14572
rect 5997 14569 6009 14572
rect 6043 14600 6055 14603
rect 8389 14603 8447 14609
rect 6043 14572 6868 14600
rect 6043 14569 6055 14572
rect 5997 14563 6055 14569
rect 1872 14532 1900 14560
rect 1872 14504 2176 14532
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14464 1639 14467
rect 1872 14464 1900 14504
rect 2038 14473 2044 14476
rect 1627 14436 1900 14464
rect 1995 14467 2044 14473
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 1995 14433 2007 14467
rect 2041 14433 2044 14467
rect 1995 14427 2044 14433
rect 2038 14424 2044 14427
rect 2096 14424 2102 14476
rect 2148 14464 2176 14504
rect 2222 14492 2228 14544
rect 2280 14532 2286 14544
rect 2869 14535 2927 14541
rect 2869 14532 2881 14535
rect 2280 14504 2881 14532
rect 2280 14492 2286 14504
rect 2869 14501 2881 14504
rect 2915 14501 2927 14535
rect 2869 14495 2927 14501
rect 4430 14492 4436 14544
rect 4488 14532 4494 14544
rect 4525 14535 4583 14541
rect 4525 14532 4537 14535
rect 4488 14504 4537 14532
rect 4488 14492 4494 14504
rect 4525 14501 4537 14504
rect 4571 14501 4583 14535
rect 4525 14495 4583 14501
rect 4614 14492 4620 14544
rect 4672 14532 4678 14544
rect 6730 14532 6736 14544
rect 4672 14504 5014 14532
rect 6691 14504 6736 14532
rect 4672 14492 4678 14504
rect 6730 14492 6736 14504
rect 6788 14492 6794 14544
rect 2593 14467 2651 14473
rect 2593 14464 2605 14467
rect 2148 14436 2605 14464
rect 2593 14433 2605 14436
rect 2639 14433 2651 14467
rect 2593 14427 2651 14433
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14433 2835 14467
rect 2958 14464 2964 14476
rect 2919 14436 2964 14464
rect 2777 14427 2835 14433
rect 1489 14399 1547 14405
rect 1489 14365 1501 14399
rect 1535 14396 1547 14399
rect 2056 14396 2084 14424
rect 2792 14396 2820 14427
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 4249 14467 4307 14473
rect 4249 14464 4261 14467
rect 4028 14436 4261 14464
rect 4028 14424 4034 14436
rect 4249 14433 4261 14436
rect 4295 14433 4307 14467
rect 4249 14427 4307 14433
rect 6457 14467 6515 14473
rect 6457 14433 6469 14467
rect 6503 14433 6515 14467
rect 6638 14464 6644 14476
rect 6599 14436 6644 14464
rect 6457 14427 6515 14433
rect 1535 14368 2820 14396
rect 1535 14365 1547 14368
rect 1489 14359 1547 14365
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 6472 14396 6500 14427
rect 6638 14424 6644 14436
rect 6696 14424 6702 14476
rect 6840 14473 6868 14572
rect 8389 14569 8401 14603
rect 8435 14600 8447 14603
rect 8938 14600 8944 14612
rect 8435 14572 8944 14600
rect 8435 14569 8447 14572
rect 8389 14563 8447 14569
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 9677 14603 9735 14609
rect 9677 14569 9689 14603
rect 9723 14600 9735 14603
rect 9766 14600 9772 14612
rect 9723 14572 9772 14600
rect 9723 14569 9735 14572
rect 9677 14563 9735 14569
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 13906 14560 13912 14612
rect 13964 14600 13970 14612
rect 14737 14603 14795 14609
rect 14737 14600 14749 14603
rect 13964 14572 14749 14600
rect 13964 14560 13970 14572
rect 14737 14569 14749 14572
rect 14783 14569 14795 14603
rect 14737 14563 14795 14569
rect 14921 14603 14979 14609
rect 14921 14569 14933 14603
rect 14967 14600 14979 14603
rect 15010 14600 15016 14612
rect 14967 14572 15016 14600
rect 14967 14569 14979 14572
rect 14921 14563 14979 14569
rect 15010 14560 15016 14572
rect 15068 14560 15074 14612
rect 7653 14535 7711 14541
rect 7653 14501 7665 14535
rect 7699 14532 7711 14535
rect 8110 14532 8116 14544
rect 7699 14504 8116 14532
rect 7699 14501 7711 14504
rect 7653 14495 7711 14501
rect 8110 14492 8116 14504
rect 8168 14532 8174 14544
rect 8481 14535 8539 14541
rect 8481 14532 8493 14535
rect 8168 14504 8493 14532
rect 8168 14492 8174 14504
rect 8481 14501 8493 14504
rect 8527 14532 8539 14535
rect 10229 14535 10287 14541
rect 10229 14532 10241 14535
rect 8527 14504 10241 14532
rect 8527 14501 8539 14504
rect 8481 14495 8539 14501
rect 10229 14501 10241 14504
rect 10275 14532 10287 14535
rect 10686 14532 10692 14544
rect 10275 14504 10692 14532
rect 10275 14501 10287 14504
rect 10229 14495 10287 14501
rect 10686 14492 10692 14504
rect 10744 14492 10750 14544
rect 12158 14492 12164 14544
rect 12216 14492 12222 14544
rect 13170 14492 13176 14544
rect 13228 14532 13234 14544
rect 13228 14504 16160 14532
rect 13228 14492 13234 14504
rect 6825 14467 6883 14473
rect 6825 14433 6837 14467
rect 6871 14433 6883 14467
rect 9490 14464 9496 14476
rect 9451 14436 9496 14464
rect 6825 14427 6883 14433
rect 9490 14424 9496 14436
rect 9548 14424 9554 14476
rect 10870 14424 10876 14476
rect 10928 14464 10934 14476
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 10928 14436 11161 14464
rect 10928 14424 10934 14436
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 11149 14427 11207 14433
rect 13817 14467 13875 14473
rect 13817 14433 13829 14467
rect 13863 14464 13875 14467
rect 14458 14464 14464 14476
rect 13863 14436 14464 14464
rect 13863 14433 13875 14436
rect 13817 14427 13875 14433
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 14918 14464 14924 14476
rect 14879 14436 14924 14464
rect 14918 14424 14924 14436
rect 14976 14464 14982 14476
rect 16132 14473 16160 14504
rect 15381 14467 15439 14473
rect 15381 14464 15393 14467
rect 14976 14436 15393 14464
rect 14976 14424 14982 14436
rect 15381 14433 15393 14436
rect 15427 14433 15439 14467
rect 15381 14427 15439 14433
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14433 16175 14467
rect 16117 14427 16175 14433
rect 5592 14368 6500 14396
rect 11425 14399 11483 14405
rect 5592 14356 5598 14368
rect 11425 14365 11437 14399
rect 11471 14396 11483 14399
rect 13078 14396 13084 14408
rect 11471 14368 13084 14396
rect 11471 14365 11483 14368
rect 11425 14359 11483 14365
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 15010 14356 15016 14408
rect 15068 14396 15074 14408
rect 15289 14399 15347 14405
rect 15289 14396 15301 14399
rect 15068 14368 15301 14396
rect 15068 14356 15074 14368
rect 15289 14365 15301 14368
rect 15335 14365 15347 14399
rect 15289 14359 15347 14365
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14365 15991 14399
rect 15933 14359 15991 14365
rect 7837 14331 7895 14337
rect 7837 14297 7849 14331
rect 7883 14328 7895 14331
rect 8938 14328 8944 14340
rect 7883 14300 8944 14328
rect 7883 14297 7895 14300
rect 7837 14291 7895 14297
rect 8938 14288 8944 14300
rect 8996 14288 9002 14340
rect 10413 14331 10471 14337
rect 10413 14297 10425 14331
rect 10459 14328 10471 14331
rect 10594 14328 10600 14340
rect 10459 14300 10600 14328
rect 10459 14297 10471 14300
rect 10413 14291 10471 14297
rect 10594 14288 10600 14300
rect 10652 14288 10658 14340
rect 12802 14288 12808 14340
rect 12860 14328 12866 14340
rect 15948 14328 15976 14359
rect 12860 14300 15976 14328
rect 12860 14288 12866 14300
rect 2133 14263 2191 14269
rect 2133 14229 2145 14263
rect 2179 14260 2191 14263
rect 5994 14260 6000 14272
rect 2179 14232 6000 14260
rect 2179 14229 2191 14232
rect 2133 14223 2191 14229
rect 5994 14220 6000 14232
rect 6052 14220 6058 14272
rect 7006 14260 7012 14272
rect 6967 14232 7012 14260
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 12894 14260 12900 14272
rect 12855 14232 12900 14260
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 13630 14260 13636 14272
rect 13591 14232 13636 14260
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 16206 14220 16212 14272
rect 16264 14260 16270 14272
rect 16301 14263 16359 14269
rect 16301 14260 16313 14263
rect 16264 14232 16313 14260
rect 16264 14220 16270 14232
rect 16301 14229 16313 14232
rect 16347 14229 16359 14263
rect 16301 14223 16359 14229
rect 1104 14170 17388 14192
rect 1104 14118 3696 14170
rect 3748 14118 3760 14170
rect 3812 14118 3824 14170
rect 3876 14118 3888 14170
rect 3940 14118 9124 14170
rect 9176 14118 9188 14170
rect 9240 14118 9252 14170
rect 9304 14118 9316 14170
rect 9368 14118 14552 14170
rect 14604 14118 14616 14170
rect 14668 14118 14680 14170
rect 14732 14118 14744 14170
rect 14796 14118 17388 14170
rect 1104 14096 17388 14118
rect 5169 14059 5227 14065
rect 5169 14025 5181 14059
rect 5215 14056 5227 14059
rect 5534 14056 5540 14068
rect 5215 14028 5540 14056
rect 5215 14025 5227 14028
rect 5169 14019 5227 14025
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 5718 14056 5724 14068
rect 5679 14028 5724 14056
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 6788 14028 6837 14056
rect 6788 14016 6794 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 6825 14019 6883 14025
rect 6932 14028 9229 14056
rect 3510 13988 3516 14000
rect 3471 13960 3516 13988
rect 3510 13948 3516 13960
rect 3568 13988 3574 14000
rect 3568 13960 4292 13988
rect 3568 13948 3574 13960
rect 4154 13920 4160 13932
rect 2884 13892 4160 13920
rect 2884 13861 2912 13892
rect 4154 13880 4160 13892
rect 4212 13880 4218 13932
rect 4264 13929 4292 13960
rect 4338 13948 4344 14000
rect 4396 13988 4402 14000
rect 6932 13988 6960 14028
rect 9217 14025 9229 14028
rect 9263 14056 9275 14059
rect 9490 14056 9496 14068
rect 9263 14028 9496 14056
rect 9263 14025 9275 14028
rect 9217 14019 9275 14025
rect 9490 14016 9496 14028
rect 9548 14056 9554 14068
rect 9769 14059 9827 14065
rect 9769 14056 9781 14059
rect 9548 14028 9781 14056
rect 9548 14016 9554 14028
rect 9769 14025 9781 14028
rect 9815 14025 9827 14059
rect 10042 14056 10048 14068
rect 10003 14028 10048 14056
rect 9769 14019 9827 14025
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 12158 14016 12164 14068
rect 12216 14056 12222 14068
rect 12253 14059 12311 14065
rect 12253 14056 12265 14059
rect 12216 14028 12265 14056
rect 12216 14016 12222 14028
rect 12253 14025 12265 14028
rect 12299 14025 12311 14059
rect 13078 14056 13084 14068
rect 13039 14028 13084 14056
rect 12253 14019 12311 14025
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 13262 14016 13268 14068
rect 13320 14056 13326 14068
rect 13633 14059 13691 14065
rect 13633 14056 13645 14059
rect 13320 14028 13645 14056
rect 13320 14016 13326 14028
rect 13633 14025 13645 14028
rect 13679 14056 13691 14059
rect 13906 14056 13912 14068
rect 13679 14028 13912 14056
rect 13679 14025 13691 14028
rect 13633 14019 13691 14025
rect 13906 14016 13912 14028
rect 13964 14016 13970 14068
rect 14366 14016 14372 14068
rect 14424 14056 14430 14068
rect 14461 14059 14519 14065
rect 14461 14056 14473 14059
rect 14424 14028 14473 14056
rect 14424 14016 14430 14028
rect 14461 14025 14473 14028
rect 14507 14025 14519 14059
rect 14461 14019 14519 14025
rect 9674 13988 9680 14000
rect 4396 13960 6960 13988
rect 8588 13960 9680 13988
rect 4396 13948 4402 13960
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 7006 13880 7012 13932
rect 7064 13920 7070 13932
rect 8588 13929 8616 13960
rect 9674 13948 9680 13960
rect 9732 13948 9738 14000
rect 13814 13988 13820 14000
rect 12452 13960 13820 13988
rect 8297 13923 8355 13929
rect 8297 13920 8309 13923
rect 7064 13892 8309 13920
rect 7064 13880 7070 13892
rect 8297 13889 8309 13892
rect 8343 13889 8355 13923
rect 8297 13883 8355 13889
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13889 8631 13923
rect 8573 13883 8631 13889
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 9640 13892 10732 13920
rect 9640 13880 9646 13892
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13821 2927 13855
rect 2869 13815 2927 13821
rect 3510 13812 3516 13864
rect 3568 13852 3574 13864
rect 3697 13855 3755 13861
rect 3697 13852 3709 13855
rect 3568 13824 3709 13852
rect 3568 13812 3574 13824
rect 3697 13821 3709 13824
rect 3743 13821 3755 13855
rect 4430 13852 4436 13864
rect 4391 13824 4436 13852
rect 3697 13815 3755 13821
rect 4430 13812 4436 13824
rect 4488 13812 4494 13864
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 5077 13855 5135 13861
rect 5077 13852 5089 13855
rect 4663 13824 5089 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 5077 13821 5089 13824
rect 5123 13852 5135 13855
rect 5596 13855 5654 13861
rect 5596 13852 5608 13855
rect 5123 13824 5608 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 5596 13821 5608 13824
rect 5642 13852 5654 13855
rect 6638 13852 6644 13864
rect 5642 13824 6644 13852
rect 5642 13821 5654 13824
rect 5596 13815 5654 13821
rect 6638 13812 6644 13824
rect 6696 13812 6702 13864
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 8938 13852 8944 13864
rect 8812 13824 8944 13852
rect 8812 13812 8818 13824
rect 8938 13812 8944 13824
rect 8996 13852 9002 13864
rect 10704 13861 10732 13892
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 8996 13824 9137 13852
rect 8996 13812 9002 13824
rect 9125 13821 9137 13824
rect 9171 13821 9183 13855
rect 9125 13815 9183 13821
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 9815 13824 9873 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 9861 13821 9873 13824
rect 9907 13821 9919 13855
rect 9861 13815 9919 13821
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13821 10747 13855
rect 11146 13852 11152 13864
rect 11107 13824 11152 13852
rect 10689 13815 10747 13821
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 12452 13861 12480 13960
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 15378 13948 15384 14000
rect 15436 13988 15442 14000
rect 15473 13991 15531 13997
rect 15473 13988 15485 13991
rect 15436 13960 15485 13988
rect 15436 13948 15442 13960
rect 15473 13957 15485 13960
rect 15519 13957 15531 13991
rect 15473 13951 15531 13957
rect 13725 13923 13783 13929
rect 13725 13920 13737 13923
rect 13556 13892 13737 13920
rect 12437 13855 12495 13861
rect 12437 13821 12449 13855
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 13262 13855 13320 13861
rect 13262 13821 13274 13855
rect 13308 13852 13320 13855
rect 13556 13852 13584 13892
rect 13725 13889 13737 13892
rect 13771 13920 13783 13923
rect 14090 13920 14096 13932
rect 13771 13892 14096 13920
rect 13771 13889 13783 13892
rect 13725 13883 13783 13889
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 13308 13824 13584 13852
rect 13308 13821 13320 13824
rect 13262 13815 13320 13821
rect 13814 13812 13820 13864
rect 13872 13852 13878 13864
rect 14277 13855 14335 13861
rect 14277 13852 14289 13855
rect 13872 13824 14289 13852
rect 13872 13812 13878 13824
rect 14277 13821 14289 13824
rect 14323 13821 14335 13855
rect 14277 13815 14335 13821
rect 15102 13812 15108 13864
rect 15160 13852 15166 13864
rect 15657 13855 15715 13861
rect 15657 13852 15669 13855
rect 15160 13824 15669 13852
rect 15160 13812 15166 13824
rect 15657 13821 15669 13824
rect 15703 13821 15715 13855
rect 16298 13852 16304 13864
rect 16259 13824 16304 13852
rect 15657 13815 15715 13821
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 7282 13744 7288 13796
rect 7340 13744 7346 13796
rect 10594 13744 10600 13796
rect 10652 13784 10658 13796
rect 13354 13784 13360 13796
rect 10652 13756 13360 13784
rect 10652 13744 10658 13756
rect 13354 13744 13360 13756
rect 13412 13744 13418 13796
rect 2682 13716 2688 13728
rect 2643 13688 2688 13716
rect 2682 13676 2688 13688
rect 2740 13676 2746 13728
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 10410 13676 10416 13728
rect 10468 13716 10474 13728
rect 10505 13719 10563 13725
rect 10505 13716 10517 13719
rect 10468 13688 10517 13716
rect 10468 13676 10474 13688
rect 10505 13685 10517 13688
rect 10551 13685 10563 13719
rect 11330 13716 11336 13728
rect 11291 13688 11336 13716
rect 10505 13679 10563 13685
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 13262 13716 13268 13728
rect 13223 13688 13268 13716
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 16022 13676 16028 13728
rect 16080 13716 16086 13728
rect 16117 13719 16175 13725
rect 16117 13716 16129 13719
rect 16080 13688 16129 13716
rect 16080 13676 16086 13688
rect 16117 13685 16129 13688
rect 16163 13685 16175 13719
rect 16117 13679 16175 13685
rect 1104 13626 17388 13648
rect 1104 13574 6410 13626
rect 6462 13574 6474 13626
rect 6526 13574 6538 13626
rect 6590 13574 6602 13626
rect 6654 13574 11838 13626
rect 11890 13574 11902 13626
rect 11954 13574 11966 13626
rect 12018 13574 12030 13626
rect 12082 13574 17388 13626
rect 1104 13552 17388 13574
rect 2958 13472 2964 13524
rect 3016 13512 3022 13524
rect 3145 13515 3203 13521
rect 3145 13512 3157 13515
rect 3016 13484 3157 13512
rect 3016 13472 3022 13484
rect 3145 13481 3157 13484
rect 3191 13481 3203 13515
rect 3145 13475 3203 13481
rect 7193 13515 7251 13521
rect 7193 13481 7205 13515
rect 7239 13512 7251 13515
rect 7282 13512 7288 13524
rect 7239 13484 7288 13512
rect 7239 13481 7251 13484
rect 7193 13475 7251 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 10042 13512 10048 13524
rect 9723 13484 10048 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 13630 13512 13636 13524
rect 10428 13484 13636 13512
rect 1394 13404 1400 13456
rect 1452 13444 1458 13456
rect 1673 13447 1731 13453
rect 1673 13444 1685 13447
rect 1452 13416 1685 13444
rect 1452 13404 1458 13416
rect 1673 13413 1685 13416
rect 1719 13413 1731 13447
rect 1673 13407 1731 13413
rect 2682 13404 2688 13456
rect 2740 13404 2746 13456
rect 4893 13447 4951 13453
rect 4893 13413 4905 13447
rect 4939 13444 4951 13447
rect 5534 13444 5540 13456
rect 4939 13416 5540 13444
rect 4939 13413 4951 13416
rect 4893 13407 4951 13413
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 10428 13444 10456 13484
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 16117 13515 16175 13521
rect 16117 13481 16129 13515
rect 16163 13512 16175 13515
rect 16482 13512 16488 13524
rect 16163 13484 16488 13512
rect 16163 13481 16175 13484
rect 16117 13475 16175 13481
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 8404 13416 10456 13444
rect 4801 13379 4859 13385
rect 4801 13345 4813 13379
rect 4847 13345 4859 13379
rect 4982 13376 4988 13388
rect 4943 13348 4988 13376
rect 4801 13339 4859 13345
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13277 1455 13311
rect 4816 13308 4844 13339
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 5166 13376 5172 13388
rect 5127 13348 5172 13376
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 6089 13379 6147 13385
rect 6089 13345 6101 13379
rect 6135 13345 6147 13379
rect 6089 13339 6147 13345
rect 7009 13379 7067 13385
rect 7009 13345 7021 13379
rect 7055 13376 7067 13379
rect 7098 13376 7104 13388
rect 7055 13348 7104 13376
rect 7055 13345 7067 13348
rect 7009 13339 7067 13345
rect 5258 13308 5264 13320
rect 4816 13280 5264 13308
rect 1397 13271 1455 13277
rect 1412 13172 1440 13271
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 6104 13308 6132 13339
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 8404 13385 8432 13416
rect 11698 13404 11704 13456
rect 11756 13404 11762 13456
rect 7837 13379 7895 13385
rect 7837 13345 7849 13379
rect 7883 13345 7895 13379
rect 7837 13339 7895 13345
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13345 8447 13379
rect 8389 13339 8447 13345
rect 9674 13379 9732 13385
rect 9674 13345 9686 13379
rect 9720 13376 9732 13379
rect 10594 13376 10600 13388
rect 9720 13348 10180 13376
rect 10555 13348 10600 13376
rect 9720 13345 9732 13348
rect 9674 13339 9732 13345
rect 7558 13308 7564 13320
rect 6104 13280 7564 13308
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 7852 13252 7880 13339
rect 10152 13320 10180 13348
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 13044 13348 13089 13376
rect 13044 13336 13050 13348
rect 13354 13336 13360 13388
rect 13412 13376 13418 13388
rect 13633 13379 13691 13385
rect 13633 13376 13645 13379
rect 13412 13348 13645 13376
rect 13412 13336 13418 13348
rect 13633 13345 13645 13348
rect 13679 13376 13691 13379
rect 14737 13379 14795 13385
rect 14737 13376 14749 13379
rect 13679 13348 14749 13376
rect 13679 13345 13691 13348
rect 13633 13339 13691 13345
rect 14737 13345 14749 13348
rect 14783 13345 14795 13379
rect 14737 13339 14795 13345
rect 16114 13379 16172 13385
rect 16114 13345 16126 13379
rect 16160 13376 16172 13379
rect 16390 13376 16396 13388
rect 16160 13348 16396 13376
rect 16160 13345 16172 13348
rect 16114 13339 16172 13345
rect 16390 13336 16396 13348
rect 16448 13376 16454 13388
rect 16577 13379 16635 13385
rect 16577 13376 16589 13379
rect 16448 13348 16589 13376
rect 16448 13336 16454 13348
rect 16577 13345 16589 13348
rect 16623 13345 16635 13379
rect 16577 13339 16635 13345
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 8205 13311 8263 13317
rect 8205 13308 8217 13311
rect 7984 13280 8217 13308
rect 7984 13268 7990 13280
rect 8205 13277 8217 13280
rect 8251 13277 8263 13311
rect 10134 13308 10140 13320
rect 10095 13280 10140 13308
rect 8205 13271 8263 13277
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 12710 13308 12716 13320
rect 12671 13280 12716 13308
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 7834 13240 7840 13252
rect 7747 13212 7840 13240
rect 7834 13200 7840 13212
rect 7892 13240 7898 13252
rect 11146 13240 11152 13252
rect 7892 13212 11152 13240
rect 7892 13200 7898 13212
rect 11146 13200 11152 13212
rect 11204 13200 11210 13252
rect 13814 13240 13820 13252
rect 13775 13212 13820 13240
rect 13814 13200 13820 13212
rect 13872 13200 13878 13252
rect 14921 13243 14979 13249
rect 14921 13209 14933 13243
rect 14967 13240 14979 13243
rect 15194 13240 15200 13252
rect 14967 13212 15200 13240
rect 14967 13209 14979 13212
rect 14921 13203 14979 13209
rect 15194 13200 15200 13212
rect 15252 13240 15258 13252
rect 16298 13240 16304 13252
rect 15252 13212 16304 13240
rect 15252 13200 15258 13212
rect 16298 13200 16304 13212
rect 16356 13200 16362 13252
rect 2958 13172 2964 13184
rect 1412 13144 2964 13172
rect 2958 13132 2964 13144
rect 3016 13132 3022 13184
rect 4617 13175 4675 13181
rect 4617 13141 4629 13175
rect 4663 13172 4675 13175
rect 4798 13172 4804 13184
rect 4663 13144 4804 13172
rect 4663 13141 4675 13144
rect 4617 13135 4675 13141
rect 4798 13132 4804 13144
rect 4856 13132 4862 13184
rect 5902 13172 5908 13184
rect 5863 13144 5908 13172
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 5994 13132 6000 13184
rect 6052 13172 6058 13184
rect 6822 13172 6828 13184
rect 6052 13144 6828 13172
rect 6052 13132 6058 13144
rect 6822 13132 6828 13144
rect 6880 13172 6886 13184
rect 7653 13175 7711 13181
rect 7653 13172 7665 13175
rect 6880 13144 7665 13172
rect 6880 13132 6886 13144
rect 7653 13141 7665 13144
rect 7699 13141 7711 13175
rect 8570 13172 8576 13184
rect 8531 13144 8576 13172
rect 7653 13135 7711 13141
rect 8570 13132 8576 13144
rect 8628 13132 8634 13184
rect 8662 13132 8668 13184
rect 8720 13172 8726 13184
rect 9490 13172 9496 13184
rect 8720 13144 9496 13172
rect 8720 13132 8726 13144
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 10042 13172 10048 13184
rect 10003 13144 10048 13172
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 10778 13172 10784 13184
rect 10739 13144 10784 13172
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 11241 13175 11299 13181
rect 11241 13141 11253 13175
rect 11287 13172 11299 13175
rect 11606 13172 11612 13184
rect 11287 13144 11612 13172
rect 11287 13141 11299 13144
rect 11241 13135 11299 13141
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 15930 13172 15936 13184
rect 15891 13144 15936 13172
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 16482 13172 16488 13184
rect 16443 13144 16488 13172
rect 16482 13132 16488 13144
rect 16540 13132 16546 13184
rect 1104 13082 17388 13104
rect 1104 13030 3696 13082
rect 3748 13030 3760 13082
rect 3812 13030 3824 13082
rect 3876 13030 3888 13082
rect 3940 13030 9124 13082
rect 9176 13030 9188 13082
rect 9240 13030 9252 13082
rect 9304 13030 9316 13082
rect 9368 13030 14552 13082
rect 14604 13030 14616 13082
rect 14668 13030 14680 13082
rect 14732 13030 14744 13082
rect 14796 13030 17388 13082
rect 1104 13008 17388 13030
rect 4614 12928 4620 12980
rect 4672 12968 4678 12980
rect 4709 12971 4767 12977
rect 4709 12968 4721 12971
rect 4672 12940 4721 12968
rect 4672 12928 4678 12940
rect 4709 12937 4721 12940
rect 4755 12968 4767 12971
rect 5166 12968 5172 12980
rect 4755 12940 5172 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 7834 12968 7840 12980
rect 7795 12940 7840 12968
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 8662 12968 8668 12980
rect 8623 12940 8668 12968
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 10134 12928 10140 12980
rect 10192 12968 10198 12980
rect 11149 12971 11207 12977
rect 11149 12968 11161 12971
rect 10192 12940 11161 12968
rect 10192 12928 10198 12940
rect 11149 12937 11161 12940
rect 11195 12937 11207 12971
rect 16390 12968 16396 12980
rect 16351 12940 16396 12968
rect 11149 12931 11207 12937
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 2317 12903 2375 12909
rect 2317 12869 2329 12903
rect 2363 12869 2375 12903
rect 2317 12863 2375 12869
rect 3605 12903 3663 12909
rect 3605 12869 3617 12903
rect 3651 12900 3663 12903
rect 4522 12900 4528 12912
rect 3651 12872 4528 12900
rect 3651 12869 3663 12872
rect 3605 12863 3663 12869
rect 1486 12832 1492 12844
rect 1447 12804 1492 12832
rect 1486 12792 1492 12804
rect 1544 12792 1550 12844
rect 1504 12696 1532 12792
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12764 1731 12767
rect 2332 12764 2360 12863
rect 4522 12860 4528 12872
rect 4580 12900 4586 12912
rect 4982 12900 4988 12912
rect 4580 12872 4988 12900
rect 4580 12860 4586 12872
rect 4982 12860 4988 12872
rect 5040 12860 5046 12912
rect 2866 12792 2872 12844
rect 2924 12832 2930 12844
rect 8757 12835 8815 12841
rect 2924 12804 3464 12832
rect 2924 12792 2930 12804
rect 1719 12736 2360 12764
rect 2501 12767 2559 12773
rect 1719 12733 1731 12736
rect 1673 12727 1731 12733
rect 2501 12733 2513 12767
rect 2547 12764 2559 12767
rect 2774 12764 2780 12776
rect 2547 12736 2780 12764
rect 2547 12733 2559 12736
rect 2501 12727 2559 12733
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 3436 12773 3464 12804
rect 5000 12804 5396 12832
rect 3329 12767 3387 12773
rect 3329 12733 3341 12767
rect 3375 12733 3387 12767
rect 3329 12727 3387 12733
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12733 3479 12767
rect 3421 12727 3479 12733
rect 3050 12696 3056 12708
rect 1504 12668 3056 12696
rect 3050 12656 3056 12668
rect 3108 12656 3114 12708
rect 3344 12696 3372 12727
rect 4154 12724 4160 12776
rect 4212 12764 4218 12776
rect 4249 12767 4307 12773
rect 4249 12764 4261 12767
rect 4212 12736 4261 12764
rect 4212 12724 4218 12736
rect 4249 12733 4261 12736
rect 4295 12733 4307 12767
rect 4249 12727 4307 12733
rect 4890 12767 4948 12773
rect 4890 12733 4902 12767
rect 4936 12764 4948 12767
rect 5000 12764 5028 12804
rect 5258 12764 5264 12776
rect 4936 12736 5028 12764
rect 5219 12736 5264 12764
rect 4936 12733 4948 12736
rect 4890 12727 4948 12733
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 5368 12773 5396 12804
rect 8757 12801 8769 12835
rect 8803 12832 8815 12835
rect 9766 12832 9772 12844
rect 8803 12804 9772 12832
rect 8803 12801 8815 12804
rect 8757 12795 8815 12801
rect 5353 12767 5411 12773
rect 5353 12733 5365 12767
rect 5399 12764 5411 12767
rect 5534 12764 5540 12776
rect 5399 12736 5540 12764
rect 5399 12733 5411 12736
rect 5353 12727 5411 12733
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 5994 12764 6000 12776
rect 5955 12736 6000 12764
rect 5994 12724 6000 12736
rect 6052 12724 6058 12776
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12733 8079 12767
rect 8021 12727 8079 12733
rect 8294 12767 8352 12773
rect 8294 12733 8306 12767
rect 8340 12764 8352 12767
rect 8570 12764 8576 12776
rect 8340 12736 8576 12764
rect 8340 12733 8352 12736
rect 8294 12727 8352 12733
rect 7282 12696 7288 12708
rect 3344 12668 7288 12696
rect 7282 12656 7288 12668
rect 7340 12696 7346 12708
rect 7926 12696 7932 12708
rect 7340 12668 7932 12696
rect 7340 12656 7346 12668
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 8036 12696 8064 12727
rect 8570 12724 8576 12736
rect 8628 12764 8634 12776
rect 8772 12764 8800 12795
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 12437 12835 12495 12841
rect 12437 12832 12449 12835
rect 10744 12804 12449 12832
rect 10744 12792 10750 12804
rect 12437 12801 12449 12804
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 14921 12835 14979 12841
rect 14921 12801 14933 12835
rect 14967 12832 14979 12835
rect 16574 12832 16580 12844
rect 14967 12804 16580 12832
rect 14967 12801 14979 12804
rect 14921 12795 14979 12801
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 9398 12764 9404 12776
rect 8628 12736 8800 12764
rect 9359 12736 9404 12764
rect 8628 12724 8634 12736
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 11330 12724 11336 12776
rect 11388 12764 11394 12776
rect 12069 12767 12127 12773
rect 12069 12764 12081 12767
rect 11388 12736 12081 12764
rect 11388 12724 11394 12736
rect 12069 12733 12081 12736
rect 12115 12733 12127 12767
rect 12069 12727 12127 12733
rect 14185 12767 14243 12773
rect 14185 12733 14197 12767
rect 14231 12764 14243 12767
rect 14645 12767 14703 12773
rect 14645 12764 14657 12767
rect 14231 12736 14657 12764
rect 14231 12733 14243 12736
rect 14185 12727 14243 12733
rect 14645 12733 14657 12736
rect 14691 12733 14703 12767
rect 14645 12727 14703 12733
rect 8478 12696 8484 12708
rect 8036 12668 8484 12696
rect 8478 12656 8484 12668
rect 8536 12656 8542 12708
rect 8662 12656 8668 12708
rect 8720 12656 8726 12708
rect 9674 12696 9680 12708
rect 9635 12668 9680 12696
rect 9674 12656 9680 12668
rect 9732 12656 9738 12708
rect 10410 12656 10416 12708
rect 10468 12656 10474 12708
rect 13630 12696 13636 12708
rect 13478 12668 13636 12696
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 13906 12696 13912 12708
rect 13867 12668 13912 12696
rect 13906 12656 13912 12668
rect 13964 12656 13970 12708
rect 1854 12628 1860 12640
rect 1815 12600 1860 12628
rect 1854 12588 1860 12600
rect 1912 12588 1918 12640
rect 4062 12628 4068 12640
rect 4023 12600 4068 12628
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 4893 12631 4951 12637
rect 4893 12597 4905 12631
rect 4939 12628 4951 12631
rect 5258 12628 5264 12640
rect 4939 12600 5264 12628
rect 4939 12597 4951 12600
rect 4893 12591 4951 12597
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5810 12628 5816 12640
rect 5771 12600 5816 12628
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8113 12631 8171 12637
rect 8113 12628 8125 12631
rect 8076 12600 8125 12628
rect 8076 12588 8082 12600
rect 8113 12597 8125 12600
rect 8159 12597 8171 12631
rect 8113 12591 8171 12597
rect 8297 12631 8355 12637
rect 8297 12597 8309 12631
rect 8343 12628 8355 12631
rect 8680 12628 8708 12656
rect 8343 12600 8708 12628
rect 8343 12597 8355 12600
rect 8297 12591 8355 12597
rect 11422 12588 11428 12640
rect 11480 12628 11486 12640
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 11480 12600 12265 12628
rect 11480 12588 11486 12600
rect 12253 12597 12265 12600
rect 12299 12628 12311 12631
rect 14200 12628 14228 12727
rect 14660 12696 14688 12727
rect 16022 12724 16028 12776
rect 16080 12724 16086 12776
rect 14918 12696 14924 12708
rect 14660 12668 14924 12696
rect 14918 12656 14924 12668
rect 14976 12656 14982 12708
rect 12299 12600 14228 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 1104 12538 17388 12560
rect 1104 12486 6410 12538
rect 6462 12486 6474 12538
rect 6526 12486 6538 12538
rect 6590 12486 6602 12538
rect 6654 12486 11838 12538
rect 11890 12486 11902 12538
rect 11954 12486 11966 12538
rect 12018 12486 12030 12538
rect 12082 12486 17388 12538
rect 1104 12464 17388 12486
rect 1394 12424 1400 12436
rect 1355 12396 1400 12424
rect 1394 12384 1400 12396
rect 1452 12384 1458 12436
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12393 1639 12427
rect 1581 12387 1639 12393
rect 1596 12356 1624 12387
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 6273 12427 6331 12433
rect 6273 12424 6285 12427
rect 5592 12396 6285 12424
rect 5592 12384 5598 12396
rect 6273 12393 6285 12396
rect 6319 12393 6331 12427
rect 6273 12387 6331 12393
rect 9582 12384 9588 12436
rect 9640 12424 9646 12436
rect 11698 12424 11704 12436
rect 9640 12396 10548 12424
rect 11659 12396 11704 12424
rect 9640 12384 9646 12396
rect 3050 12356 3056 12368
rect 1596 12328 1992 12356
rect 3011 12328 3056 12356
rect 1578 12291 1636 12297
rect 1578 12257 1590 12291
rect 1624 12288 1636 12291
rect 1854 12288 1860 12300
rect 1624 12260 1860 12288
rect 1624 12257 1636 12260
rect 1578 12251 1636 12257
rect 1854 12248 1860 12260
rect 1912 12248 1918 12300
rect 1964 12297 1992 12328
rect 3050 12316 3056 12328
rect 3108 12316 3114 12368
rect 4798 12356 4804 12368
rect 4759 12328 4804 12356
rect 4798 12316 4804 12328
rect 4856 12316 4862 12368
rect 6914 12316 6920 12368
rect 6972 12356 6978 12368
rect 7009 12359 7067 12365
rect 7009 12356 7021 12359
rect 6972 12328 7021 12356
rect 6972 12316 6978 12328
rect 7009 12325 7021 12328
rect 7055 12325 7067 12359
rect 7009 12319 7067 12325
rect 7742 12316 7748 12368
rect 7800 12316 7806 12368
rect 9677 12359 9735 12365
rect 9677 12325 9689 12359
rect 9723 12356 9735 12359
rect 9950 12356 9956 12368
rect 9723 12328 9956 12356
rect 9723 12325 9735 12328
rect 9677 12319 9735 12325
rect 9950 12316 9956 12328
rect 10008 12316 10014 12368
rect 10520 12365 10548 12396
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 12345 12427 12403 12433
rect 12345 12393 12357 12427
rect 12391 12424 12403 12427
rect 12434 12424 12440 12436
rect 12391 12396 12440 12424
rect 12391 12393 12403 12396
rect 12345 12387 12403 12393
rect 12434 12384 12440 12396
rect 12492 12424 12498 12436
rect 12894 12424 12900 12436
rect 12492 12396 12900 12424
rect 12492 12384 12498 12396
rect 10505 12359 10563 12365
rect 10505 12325 10517 12359
rect 10551 12325 10563 12359
rect 10505 12319 10563 12325
rect 10594 12316 10600 12368
rect 10652 12356 10658 12368
rect 10689 12359 10747 12365
rect 10689 12356 10701 12359
rect 10652 12328 10701 12356
rect 10652 12316 10658 12328
rect 10689 12325 10701 12328
rect 10735 12325 10747 12359
rect 10689 12319 10747 12325
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2130 12288 2136 12300
rect 1995 12260 2136 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 3237 12291 3295 12297
rect 3237 12257 3249 12291
rect 3283 12288 3295 12291
rect 3510 12288 3516 12300
rect 3283 12260 3516 12288
rect 3283 12257 3295 12260
rect 3237 12251 3295 12257
rect 3510 12248 3516 12260
rect 3568 12248 3574 12300
rect 5902 12248 5908 12300
rect 5960 12248 5966 12300
rect 9490 12288 9496 12300
rect 9451 12260 9496 12288
rect 9490 12248 9496 12260
rect 9548 12248 9554 12300
rect 9769 12291 9827 12297
rect 9769 12257 9781 12291
rect 9815 12257 9827 12291
rect 9769 12251 9827 12257
rect 1872 12220 1900 12248
rect 2041 12223 2099 12229
rect 2041 12220 2053 12223
rect 1872 12192 2053 12220
rect 2041 12189 2053 12192
rect 2087 12220 2099 12223
rect 2222 12220 2228 12232
rect 2087 12192 2228 12220
rect 2087 12189 2099 12192
rect 2041 12183 2099 12189
rect 2222 12180 2228 12192
rect 2280 12180 2286 12232
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 3016 12192 4537 12220
rect 3016 12180 3022 12192
rect 4525 12189 4537 12192
rect 4571 12220 4583 12223
rect 5534 12220 5540 12232
rect 4571 12192 5540 12220
rect 4571 12189 4583 12192
rect 4525 12183 4583 12189
rect 5534 12180 5540 12192
rect 5592 12220 5598 12232
rect 5810 12220 5816 12232
rect 5592 12192 5816 12220
rect 5592 12180 5598 12192
rect 5810 12180 5816 12192
rect 5868 12220 5874 12232
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 5868 12192 6745 12220
rect 5868 12180 5874 12192
rect 6733 12189 6745 12192
rect 6779 12189 6791 12223
rect 9784 12220 9812 12251
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 11517 12291 11575 12297
rect 9916 12260 9961 12288
rect 9916 12248 9922 12260
rect 11517 12257 11529 12291
rect 11563 12257 11575 12291
rect 11517 12251 11575 12257
rect 10134 12220 10140 12232
rect 9784 12192 10140 12220
rect 6733 12183 6791 12189
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 10045 12155 10103 12161
rect 10045 12152 10057 12155
rect 9732 12124 10057 12152
rect 9732 12112 9738 12124
rect 10045 12121 10057 12124
rect 10091 12121 10103 12155
rect 11532 12152 11560 12251
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 12342 12297 12348 12300
rect 12286 12291 12348 12297
rect 12286 12288 12298 12291
rect 11664 12260 12298 12288
rect 11664 12248 11670 12260
rect 12286 12257 12298 12260
rect 12332 12257 12348 12291
rect 12286 12251 12348 12257
rect 12342 12248 12348 12251
rect 12400 12248 12406 12300
rect 12728 12297 12756 12396
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 13630 12424 13636 12436
rect 13591 12396 13636 12424
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 13906 12384 13912 12436
rect 13964 12424 13970 12436
rect 14921 12427 14979 12433
rect 14921 12424 14933 12427
rect 13964 12396 14933 12424
rect 13964 12384 13970 12396
rect 14921 12393 14933 12396
rect 14967 12393 14979 12427
rect 14921 12387 14979 12393
rect 15105 12427 15163 12433
rect 15105 12393 15117 12427
rect 15151 12424 15163 12427
rect 15151 12396 15516 12424
rect 15151 12393 15163 12396
rect 15105 12387 15163 12393
rect 15194 12356 15200 12368
rect 13832 12328 15200 12356
rect 13832 12297 13860 12328
rect 15194 12316 15200 12328
rect 15252 12316 15258 12368
rect 15488 12297 15516 12396
rect 16390 12384 16396 12436
rect 16448 12384 16454 12436
rect 16574 12424 16580 12436
rect 16535 12396 16580 12424
rect 16574 12384 16580 12396
rect 16632 12384 16638 12436
rect 16206 12356 16212 12368
rect 16167 12328 16212 12356
rect 16206 12316 16212 12328
rect 16264 12316 16270 12368
rect 16301 12359 16359 12365
rect 16301 12325 16313 12359
rect 16347 12356 16359 12359
rect 16408 12356 16436 12384
rect 16347 12328 16436 12356
rect 16347 12325 16359 12328
rect 16301 12319 16359 12325
rect 12713 12291 12771 12297
rect 12713 12257 12725 12291
rect 12759 12257 12771 12291
rect 12713 12251 12771 12257
rect 13817 12291 13875 12297
rect 13817 12257 13829 12291
rect 13863 12257 13875 12291
rect 13817 12251 13875 12257
rect 15102 12291 15160 12297
rect 15102 12257 15114 12291
rect 15148 12288 15160 12291
rect 15473 12291 15531 12297
rect 15148 12260 15424 12288
rect 15148 12257 15160 12260
rect 15102 12251 15160 12257
rect 12357 12220 12385 12248
rect 12805 12223 12863 12229
rect 12805 12220 12817 12223
rect 12357 12192 12817 12220
rect 12805 12189 12817 12192
rect 12851 12189 12863 12223
rect 15396 12220 15424 12260
rect 15473 12257 15485 12291
rect 15519 12288 15531 12291
rect 15930 12288 15936 12300
rect 15519 12260 15936 12288
rect 15519 12257 15531 12260
rect 15473 12251 15531 12257
rect 15930 12248 15936 12260
rect 15988 12288 15994 12300
rect 16025 12291 16083 12297
rect 16025 12288 16037 12291
rect 15988 12260 16037 12288
rect 15988 12248 15994 12260
rect 16025 12257 16037 12260
rect 16071 12257 16083 12291
rect 16025 12251 16083 12257
rect 15565 12223 15623 12229
rect 15565 12220 15577 12223
rect 15396 12192 15577 12220
rect 12805 12183 12863 12189
rect 15565 12189 15577 12192
rect 15611 12220 15623 12223
rect 16224 12220 16252 12316
rect 16393 12291 16451 12297
rect 16393 12257 16405 12291
rect 16439 12288 16451 12291
rect 16482 12288 16488 12300
rect 16439 12260 16488 12288
rect 16439 12257 16451 12260
rect 16393 12251 16451 12257
rect 16482 12248 16488 12260
rect 16540 12248 16546 12300
rect 15611 12192 16252 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 11532 12124 12434 12152
rect 10045 12115 10103 12121
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 4338 12084 4344 12096
rect 3568 12056 4344 12084
rect 3568 12044 3574 12056
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 8481 12087 8539 12093
rect 8481 12053 8493 12087
rect 8527 12084 8539 12087
rect 9858 12084 9864 12096
rect 8527 12056 9864 12084
rect 8527 12053 8539 12056
rect 8481 12047 8539 12053
rect 9858 12044 9864 12056
rect 9916 12044 9922 12096
rect 12066 12044 12072 12096
rect 12124 12084 12130 12096
rect 12161 12087 12219 12093
rect 12161 12084 12173 12087
rect 12124 12056 12173 12084
rect 12124 12044 12130 12056
rect 12161 12053 12173 12056
rect 12207 12053 12219 12087
rect 12406 12084 12434 12124
rect 13354 12084 13360 12096
rect 12406 12056 13360 12084
rect 12161 12047 12219 12053
rect 13354 12044 13360 12056
rect 13412 12084 13418 12096
rect 13814 12084 13820 12096
rect 13412 12056 13820 12084
rect 13412 12044 13418 12056
rect 13814 12044 13820 12056
rect 13872 12044 13878 12096
rect 1104 11994 17388 12016
rect 1104 11942 3696 11994
rect 3748 11942 3760 11994
rect 3812 11942 3824 11994
rect 3876 11942 3888 11994
rect 3940 11942 9124 11994
rect 9176 11942 9188 11994
rect 9240 11942 9252 11994
rect 9304 11942 9316 11994
rect 9368 11942 14552 11994
rect 14604 11942 14616 11994
rect 14668 11942 14680 11994
rect 14732 11942 14744 11994
rect 14796 11942 17388 11994
rect 1104 11920 17388 11942
rect 4614 11880 4620 11892
rect 4575 11852 4620 11880
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 7742 11880 7748 11892
rect 7703 11852 7748 11880
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 10597 11883 10655 11889
rect 10597 11849 10609 11883
rect 10643 11880 10655 11883
rect 10686 11880 10692 11892
rect 10643 11852 10692 11880
rect 10643 11849 10655 11852
rect 10597 11843 10655 11849
rect 10686 11840 10692 11852
rect 10744 11840 10750 11892
rect 12621 11883 12679 11889
rect 12621 11849 12633 11883
rect 12667 11880 12679 11883
rect 12710 11880 12716 11892
rect 12667 11852 12716 11880
rect 12667 11849 12679 11852
rect 12621 11843 12679 11849
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11744 2375 11747
rect 2958 11744 2964 11756
rect 2363 11716 2964 11744
rect 2363 11713 2375 11716
rect 2317 11707 2375 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 4522 11744 4528 11756
rect 4483 11716 4528 11744
rect 4522 11704 4528 11716
rect 4580 11704 4586 11756
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 11422 11744 11428 11756
rect 9548 11716 11428 11744
rect 9548 11704 9554 11716
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 14918 11704 14924 11756
rect 14976 11744 14982 11756
rect 15749 11747 15807 11753
rect 15749 11744 15761 11747
rect 14976 11716 15761 11744
rect 14976 11704 14982 11716
rect 15749 11713 15761 11716
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 4062 11676 4068 11688
rect 3726 11648 4068 11676
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4540 11676 4568 11704
rect 4988 11679 5046 11685
rect 4988 11676 5000 11679
rect 4540 11648 5000 11676
rect 4988 11645 5000 11648
rect 5034 11645 5046 11679
rect 7558 11676 7564 11688
rect 7519 11648 7564 11676
rect 4988 11639 5046 11645
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 10226 11679 10284 11685
rect 10226 11645 10238 11679
rect 10272 11676 10284 11679
rect 10594 11676 10600 11688
rect 10272 11648 10600 11676
rect 10272 11645 10284 11648
rect 10226 11639 10284 11645
rect 10594 11636 10600 11648
rect 10652 11676 10658 11688
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 10652 11648 10701 11676
rect 10652 11636 10658 11648
rect 10689 11645 10701 11648
rect 10735 11645 10747 11679
rect 12066 11676 12072 11688
rect 12027 11648 12072 11676
rect 10689 11639 10747 11645
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 12342 11676 12348 11688
rect 12303 11648 12348 11676
rect 12342 11636 12348 11648
rect 12400 11636 12406 11688
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 16390 11676 16396 11688
rect 12492 11648 12537 11676
rect 16351 11648 16396 11676
rect 12492 11636 12498 11648
rect 16390 11636 16396 11648
rect 16448 11636 16454 11688
rect 2590 11608 2596 11620
rect 2551 11580 2596 11608
rect 2590 11568 2596 11580
rect 2648 11568 2654 11620
rect 12250 11608 12256 11620
rect 12211 11580 12256 11608
rect 12250 11568 12256 11580
rect 12308 11568 12314 11620
rect 13814 11568 13820 11620
rect 13872 11608 13878 11620
rect 15470 11608 15476 11620
rect 13872 11580 14306 11608
rect 15431 11580 15476 11608
rect 13872 11568 13878 11580
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 2682 11500 2688 11552
rect 2740 11540 2746 11552
rect 4065 11543 4123 11549
rect 4065 11540 4077 11543
rect 2740 11512 4077 11540
rect 2740 11500 2746 11512
rect 4065 11509 4077 11512
rect 4111 11509 4123 11543
rect 4065 11503 4123 11509
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 4985 11543 5043 11549
rect 4985 11540 4997 11543
rect 4672 11512 4997 11540
rect 4672 11500 4678 11512
rect 4985 11509 4997 11512
rect 5031 11509 5043 11543
rect 4985 11503 5043 11509
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5169 11543 5227 11549
rect 5169 11540 5181 11543
rect 5132 11512 5181 11540
rect 5132 11500 5138 11512
rect 5169 11509 5181 11512
rect 5215 11509 5227 11543
rect 10042 11540 10048 11552
rect 10003 11512 10048 11540
rect 5169 11503 5227 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10229 11543 10287 11549
rect 10229 11509 10241 11543
rect 10275 11540 10287 11543
rect 10686 11540 10692 11552
rect 10275 11512 10692 11540
rect 10275 11509 10287 11512
rect 10229 11503 10287 11509
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 13998 11540 14004 11552
rect 13959 11512 14004 11540
rect 13998 11500 14004 11512
rect 14056 11500 14062 11552
rect 16206 11540 16212 11552
rect 16167 11512 16212 11540
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 1104 11450 17388 11472
rect 1104 11398 6410 11450
rect 6462 11398 6474 11450
rect 6526 11398 6538 11450
rect 6590 11398 6602 11450
rect 6654 11398 11838 11450
rect 11890 11398 11902 11450
rect 11954 11398 11966 11450
rect 12018 11398 12030 11450
rect 12082 11398 17388 11450
rect 1104 11376 17388 11398
rect 2130 11336 2136 11348
rect 2091 11308 2136 11336
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2406 11336 2412 11348
rect 2363 11308 2412 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 5626 11336 5632 11348
rect 3988 11308 5632 11336
rect 1762 11200 1768 11212
rect 1723 11172 1768 11200
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 2314 11200 2320 11212
rect 2227 11172 2320 11200
rect 2314 11160 2320 11172
rect 2372 11200 2378 11212
rect 2682 11200 2688 11212
rect 2372 11172 2688 11200
rect 2372 11160 2378 11172
rect 2682 11160 2688 11172
rect 2740 11200 2746 11212
rect 2777 11203 2835 11209
rect 2777 11200 2789 11203
rect 2740 11172 2789 11200
rect 2740 11160 2746 11172
rect 2777 11169 2789 11172
rect 2823 11169 2835 11203
rect 2777 11163 2835 11169
rect 3988 11132 4016 11308
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 6273 11339 6331 11345
rect 6273 11305 6285 11339
rect 6319 11336 6331 11339
rect 7101 11339 7159 11345
rect 7101 11336 7113 11339
rect 6319 11308 7113 11336
rect 6319 11305 6331 11308
rect 6273 11299 6331 11305
rect 7101 11305 7113 11308
rect 7147 11336 7159 11339
rect 7466 11336 7472 11348
rect 7147 11308 7472 11336
rect 7147 11305 7159 11308
rect 7101 11299 7159 11305
rect 7466 11296 7472 11308
rect 7524 11296 7530 11348
rect 12158 11296 12164 11348
rect 12216 11336 12222 11348
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 12216 11308 12265 11336
rect 12216 11296 12222 11308
rect 12253 11305 12265 11308
rect 12299 11305 12311 11339
rect 13814 11336 13820 11348
rect 13775 11308 13820 11336
rect 12253 11299 12311 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 16540 11308 16681 11336
rect 16540 11296 16546 11308
rect 16669 11305 16681 11308
rect 16715 11305 16727 11339
rect 16669 11299 16727 11305
rect 4801 11271 4859 11277
rect 4801 11237 4813 11271
rect 4847 11268 4859 11271
rect 5074 11268 5080 11280
rect 4847 11240 5080 11268
rect 4847 11237 4859 11240
rect 4801 11231 4859 11237
rect 5074 11228 5080 11240
rect 5132 11228 5138 11280
rect 5810 11228 5816 11280
rect 5868 11228 5874 11280
rect 9582 11228 9588 11280
rect 9640 11228 9646 11280
rect 11330 11268 11336 11280
rect 10626 11240 11336 11268
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 7098 11203 7156 11209
rect 7098 11169 7110 11203
rect 7144 11200 7156 11203
rect 8570 11200 8576 11212
rect 7144 11172 7420 11200
rect 8483 11172 8576 11200
rect 7144 11169 7156 11172
rect 7098 11163 7156 11169
rect 7392 11144 7420 11172
rect 8570 11160 8576 11172
rect 8628 11200 8634 11212
rect 9600 11200 9628 11228
rect 8628 11172 9628 11200
rect 11885 11203 11943 11209
rect 8628 11160 8634 11172
rect 11885 11169 11897 11203
rect 11931 11200 11943 11203
rect 12176 11200 12204 11296
rect 15194 11268 15200 11280
rect 13648 11240 15200 11268
rect 11931 11172 12204 11200
rect 11931 11169 11943 11172
rect 11885 11163 11943 11169
rect 12250 11160 12256 11212
rect 12308 11200 12314 11212
rect 12897 11203 12955 11209
rect 12308 11172 12401 11200
rect 12308 11160 12314 11172
rect 12897 11169 12909 11203
rect 12943 11200 12955 11203
rect 13354 11200 13360 11212
rect 12943 11172 13360 11200
rect 12943 11169 12955 11172
rect 12897 11163 12955 11169
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 13648 11209 13676 11240
rect 15194 11228 15200 11240
rect 15252 11228 15258 11280
rect 16206 11228 16212 11280
rect 16264 11228 16270 11280
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11169 13691 11203
rect 14918 11200 14924 11212
rect 14879 11172 14924 11200
rect 13633 11163 13691 11169
rect 14918 11160 14924 11172
rect 14976 11160 14982 11212
rect 1964 11104 4016 11132
rect 1964 11073 1992 11104
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 4120 11104 4537 11132
rect 4120 11092 4126 11104
rect 4525 11101 4537 11104
rect 4571 11132 4583 11135
rect 5534 11132 5540 11144
rect 4571 11104 5540 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7432 11104 7573 11132
rect 7432 11092 7438 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11132 9643 11135
rect 10594 11132 10600 11144
rect 9631 11104 10600 11132
rect 9631 11101 9643 11104
rect 9585 11095 9643 11101
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 11054 11132 11060 11144
rect 11015 11104 11060 11132
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11132 11391 11135
rect 11422 11132 11428 11144
rect 11379 11104 11428 11132
rect 11379 11101 11391 11104
rect 11333 11095 11391 11101
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 11698 11092 11704 11144
rect 11756 11132 11762 11144
rect 11793 11135 11851 11141
rect 11793 11132 11805 11135
rect 11756 11104 11805 11132
rect 11756 11092 11762 11104
rect 11793 11101 11805 11104
rect 11839 11132 11851 11135
rect 12268 11132 12296 11160
rect 11839 11104 12296 11132
rect 11839 11101 11851 11104
rect 11793 11095 11851 11101
rect 1949 11067 2007 11073
rect 1949 11033 1961 11067
rect 1995 11033 2007 11067
rect 7466 11064 7472 11076
rect 7427 11036 7472 11064
rect 1949 11027 2007 11033
rect 7466 11024 7472 11036
rect 7524 11024 7530 11076
rect 8386 11064 8392 11076
rect 8347 11036 8392 11064
rect 8386 11024 8392 11036
rect 8444 11024 8450 11076
rect 13078 11064 13084 11076
rect 13039 11036 13084 11064
rect 13078 11024 13084 11036
rect 13136 11024 13142 11076
rect 2406 10956 2412 11008
rect 2464 10996 2470 11008
rect 2685 10999 2743 11005
rect 2685 10996 2697 10999
rect 2464 10968 2697 10996
rect 2464 10956 2470 10968
rect 2685 10965 2697 10968
rect 2731 10965 2743 10999
rect 2685 10959 2743 10965
rect 6917 10999 6975 11005
rect 6917 10965 6929 10999
rect 6963 10996 6975 10999
rect 7006 10996 7012 11008
rect 6963 10968 7012 10996
rect 6963 10965 6975 10968
rect 6917 10959 6975 10965
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 7558 10996 7564 11008
rect 7156 10968 7564 10996
rect 7156 10956 7162 10968
rect 7558 10956 7564 10968
rect 7616 10996 7622 11008
rect 10870 10996 10876 11008
rect 7616 10968 10876 10996
rect 7616 10956 7622 10968
rect 10870 10956 10876 10968
rect 10928 10956 10934 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 15194 11005 15200 11008
rect 15184 10999 15200 11005
rect 12492 10968 12537 10996
rect 12492 10956 12498 10968
rect 15184 10965 15196 10999
rect 15184 10959 15200 10965
rect 15194 10956 15200 10959
rect 15252 10956 15258 11008
rect 1104 10906 17388 10928
rect 1104 10854 3696 10906
rect 3748 10854 3760 10906
rect 3812 10854 3824 10906
rect 3876 10854 3888 10906
rect 3940 10854 9124 10906
rect 9176 10854 9188 10906
rect 9240 10854 9252 10906
rect 9304 10854 9316 10906
rect 9368 10854 14552 10906
rect 14604 10854 14616 10906
rect 14668 10854 14680 10906
rect 14732 10854 14744 10906
rect 14796 10854 17388 10906
rect 1104 10832 17388 10854
rect 2590 10792 2596 10804
rect 2551 10764 2596 10792
rect 2590 10752 2596 10764
rect 2648 10752 2654 10804
rect 4062 10792 4068 10804
rect 3712 10764 4068 10792
rect 3712 10665 3740 10764
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 5258 10752 5264 10804
rect 5316 10792 5322 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 5316 10764 5457 10792
rect 5316 10752 5322 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 10100 10764 10149 10792
rect 10100 10752 10106 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 10137 10755 10195 10761
rect 10873 10795 10931 10801
rect 10873 10761 10885 10795
rect 10919 10792 10931 10795
rect 11054 10792 11060 10804
rect 10919 10764 11060 10792
rect 10919 10761 10931 10764
rect 10873 10755 10931 10761
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11330 10792 11336 10804
rect 11291 10764 11336 10792
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 15381 10795 15439 10801
rect 15381 10761 15393 10795
rect 15427 10792 15439 10795
rect 15470 10792 15476 10804
rect 15427 10764 15476 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 9585 10727 9643 10733
rect 9585 10693 9597 10727
rect 9631 10693 9643 10727
rect 9585 10687 9643 10693
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10656 4031 10659
rect 9600 10656 9628 10687
rect 13630 10684 13636 10736
rect 13688 10724 13694 10736
rect 13688 10696 15792 10724
rect 13688 10684 13694 10696
rect 4019 10628 9628 10656
rect 10244 10628 10548 10656
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 2130 10588 2136 10600
rect 2087 10560 2136 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2130 10548 2136 10560
rect 2188 10548 2194 10600
rect 2222 10548 2228 10600
rect 2280 10588 2286 10600
rect 2406 10588 2412 10600
rect 2280 10560 2325 10588
rect 2367 10560 2412 10588
rect 2280 10548 2286 10560
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 3234 10588 3240 10600
rect 3195 10560 3240 10588
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 5074 10548 5080 10600
rect 5132 10548 5138 10600
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 9490 10588 9496 10600
rect 9171 10560 9496 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 9674 10548 9680 10600
rect 9732 10597 9738 10600
rect 10244 10597 10272 10628
rect 10520 10597 10548 10628
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 12069 10659 12127 10665
rect 12069 10656 12081 10659
rect 11480 10628 12081 10656
rect 11480 10616 11486 10628
rect 12069 10625 12081 10628
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 12345 10659 12403 10665
rect 12345 10625 12357 10659
rect 12391 10656 12403 10659
rect 12434 10656 12440 10668
rect 12391 10628 12440 10656
rect 12391 10625 12403 10628
rect 12345 10619 12403 10625
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10656 13875 10659
rect 14369 10659 14427 10665
rect 14369 10656 14381 10659
rect 13863 10628 14381 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 9732 10591 9768 10597
rect 9756 10588 9768 10591
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 9756 10560 10241 10588
rect 9756 10557 9768 10560
rect 9732 10551 9768 10557
rect 10229 10557 10241 10560
rect 10275 10557 10287 10591
rect 10229 10551 10287 10557
rect 10321 10591 10379 10597
rect 10321 10557 10333 10591
rect 10367 10557 10379 10591
rect 10321 10551 10379 10557
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10557 10563 10591
rect 10686 10588 10692 10600
rect 10647 10560 10692 10588
rect 10505 10551 10563 10557
rect 9732 10548 9738 10551
rect 2314 10520 2320 10532
rect 2275 10492 2320 10520
rect 2314 10480 2320 10492
rect 2372 10480 2378 10532
rect 8386 10480 8392 10532
rect 8444 10480 8450 10532
rect 8846 10520 8852 10532
rect 8807 10492 8852 10520
rect 8846 10480 8852 10492
rect 8904 10480 8910 10532
rect 10042 10520 10048 10532
rect 9784 10492 10048 10520
rect 3050 10452 3056 10464
rect 3011 10424 3056 10452
rect 3050 10412 3056 10424
rect 3108 10412 3114 10464
rect 7374 10452 7380 10464
rect 7335 10424 7380 10452
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 9784 10461 9812 10492
rect 10042 10480 10048 10492
rect 10100 10520 10106 10532
rect 10336 10520 10364 10551
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 10778 10548 10784 10600
rect 10836 10588 10842 10600
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 10836 10560 11529 10588
rect 10836 10548 10842 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 10100 10492 10364 10520
rect 10100 10480 10106 10492
rect 10594 10480 10600 10532
rect 10652 10520 10658 10532
rect 10652 10492 10697 10520
rect 10652 10480 10658 10492
rect 13078 10480 13084 10532
rect 13136 10480 13142 10532
rect 9769 10455 9827 10461
rect 9769 10421 9781 10455
rect 9815 10421 9827 10455
rect 13924 10452 13952 10628
rect 14369 10625 14381 10628
rect 14415 10625 14427 10659
rect 14369 10619 14427 10625
rect 15304 10628 15700 10656
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 14056 10560 14289 10588
rect 14056 10548 14062 10560
rect 14277 10557 14289 10560
rect 14323 10588 14335 10591
rect 14740 10591 14798 10597
rect 14740 10588 14752 10591
rect 14323 10560 14752 10588
rect 14323 10557 14335 10560
rect 14277 10551 14335 10557
rect 14740 10557 14752 10560
rect 14786 10588 14798 10591
rect 15304 10588 15332 10628
rect 15672 10597 15700 10628
rect 15764 10597 15792 10696
rect 14786 10560 15332 10588
rect 15565 10591 15623 10597
rect 14786 10557 14798 10560
rect 14740 10551 14798 10557
rect 15565 10557 15577 10591
rect 15611 10557 15623 10591
rect 15565 10551 15623 10557
rect 15657 10591 15715 10597
rect 15657 10557 15669 10591
rect 15703 10557 15715 10591
rect 15657 10551 15715 10557
rect 15749 10591 15807 10597
rect 15749 10557 15761 10591
rect 15795 10557 15807 10591
rect 15749 10551 15807 10557
rect 15933 10591 15991 10597
rect 15933 10557 15945 10591
rect 15979 10557 15991 10591
rect 15933 10551 15991 10557
rect 15580 10520 15608 10551
rect 14752 10492 15608 10520
rect 14752 10461 14780 10492
rect 14737 10455 14795 10461
rect 14737 10452 14749 10455
rect 13924 10424 14749 10452
rect 9769 10415 9827 10421
rect 14737 10421 14749 10424
rect 14783 10421 14795 10455
rect 14918 10452 14924 10464
rect 14831 10424 14924 10452
rect 14737 10415 14795 10421
rect 14918 10412 14924 10424
rect 14976 10452 14982 10464
rect 15948 10452 15976 10551
rect 14976 10424 15976 10452
rect 14976 10412 14982 10424
rect 1104 10362 17388 10384
rect 1104 10310 6410 10362
rect 6462 10310 6474 10362
rect 6526 10310 6538 10362
rect 6590 10310 6602 10362
rect 6654 10310 11838 10362
rect 11890 10310 11902 10362
rect 11954 10310 11966 10362
rect 12018 10310 12030 10362
rect 12082 10310 17388 10362
rect 1104 10288 17388 10310
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10248 3203 10251
rect 3326 10248 3332 10260
rect 3191 10220 3332 10248
rect 3191 10217 3203 10220
rect 3145 10211 3203 10217
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 5074 10208 5080 10260
rect 5132 10248 5138 10260
rect 5169 10251 5227 10257
rect 5169 10248 5181 10251
rect 5132 10220 5181 10248
rect 5132 10208 5138 10220
rect 5169 10217 5181 10220
rect 5215 10217 5227 10251
rect 5810 10248 5816 10260
rect 5771 10220 5816 10248
rect 5169 10211 5227 10217
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 6825 10251 6883 10257
rect 6825 10217 6837 10251
rect 6871 10248 6883 10251
rect 6914 10248 6920 10260
rect 6871 10220 6920 10248
rect 6871 10217 6883 10220
rect 6825 10211 6883 10217
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7064 10220 7328 10248
rect 7064 10208 7070 10220
rect 1394 10140 1400 10192
rect 1452 10180 1458 10192
rect 1673 10183 1731 10189
rect 1673 10180 1685 10183
rect 1452 10152 1685 10180
rect 1452 10140 1458 10152
rect 1673 10149 1685 10152
rect 1719 10149 1731 10183
rect 3050 10180 3056 10192
rect 2898 10152 3056 10180
rect 1673 10143 1731 10149
rect 3050 10140 3056 10152
rect 3108 10140 3114 10192
rect 7098 10180 7104 10192
rect 6012 10152 7104 10180
rect 6012 10121 6040 10152
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 5997 10115 6055 10121
rect 5997 10112 6009 10115
rect 5399 10084 6009 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 5997 10081 6009 10084
rect 6043 10081 6055 10115
rect 5997 10075 6055 10081
rect 7006 10115 7064 10121
rect 7006 10081 7018 10115
rect 7052 10112 7064 10115
rect 7300 10112 7328 10220
rect 7466 10208 7472 10260
rect 7524 10248 7530 10260
rect 8481 10251 8539 10257
rect 7524 10220 8340 10248
rect 7524 10208 7530 10220
rect 7374 10140 7380 10192
rect 7432 10180 7438 10192
rect 8205 10183 8263 10189
rect 8205 10180 8217 10183
rect 7432 10152 8217 10180
rect 7432 10140 7438 10152
rect 8205 10149 8217 10152
rect 8251 10149 8263 10183
rect 8205 10143 8263 10149
rect 7929 10115 7987 10121
rect 7929 10112 7941 10115
rect 7052 10084 7236 10112
rect 7052 10081 7064 10084
rect 7006 10075 7064 10081
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 2958 10044 2964 10056
rect 1443 10016 2964 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 7208 9976 7236 10084
rect 7300 10084 7941 10112
rect 7300 10044 7328 10084
rect 7929 10081 7941 10084
rect 7975 10081 7987 10115
rect 8110 10112 8116 10124
rect 8071 10084 8116 10112
rect 7929 10075 7987 10081
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 8312 10121 8340 10220
rect 8481 10217 8493 10251
rect 8527 10248 8539 10251
rect 8846 10248 8852 10260
rect 8527 10220 8852 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 11698 10248 11704 10260
rect 11659 10220 11704 10248
rect 11698 10208 11704 10220
rect 11756 10208 11762 10260
rect 13173 10251 13231 10257
rect 13173 10217 13185 10251
rect 13219 10248 13231 10251
rect 13219 10220 13584 10248
rect 13219 10217 13231 10220
rect 13173 10211 13231 10217
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10081 8355 10115
rect 8297 10075 8355 10081
rect 8938 10072 8944 10124
rect 8996 10112 9002 10124
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 8996 10084 9505 10112
rect 8996 10072 9002 10084
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 11146 10072 11152 10124
rect 11204 10112 11210 10124
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 11204 10084 11897 10112
rect 11204 10072 11210 10084
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 11885 10075 11943 10081
rect 12069 10115 12127 10121
rect 12069 10081 12081 10115
rect 12115 10112 12127 10115
rect 12802 10112 12808 10124
rect 12115 10084 12808 10112
rect 12115 10081 12127 10084
rect 12069 10075 12127 10081
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 13170 10112 13176 10124
rect 13083 10084 13176 10112
rect 13170 10072 13176 10084
rect 13228 10112 13234 10124
rect 13556 10121 13584 10220
rect 15657 10183 15715 10189
rect 15657 10149 15669 10183
rect 15703 10180 15715 10183
rect 15746 10180 15752 10192
rect 15703 10152 15752 10180
rect 15703 10149 15715 10152
rect 15657 10143 15715 10149
rect 15746 10140 15752 10152
rect 15804 10140 15810 10192
rect 13541 10115 13599 10121
rect 13228 10084 13492 10112
rect 13228 10072 13234 10084
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 7300 10016 7389 10044
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7377 10007 7435 10013
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10044 7527 10047
rect 8128 10044 8156 10072
rect 7515 10016 8156 10044
rect 13464 10044 13492 10084
rect 13541 10081 13553 10115
rect 13587 10112 13599 10115
rect 14918 10112 14924 10124
rect 13587 10084 14924 10112
rect 13587 10081 13599 10084
rect 13541 10075 13599 10081
rect 14918 10072 14924 10084
rect 14976 10072 14982 10124
rect 15470 10112 15476 10124
rect 15431 10084 15476 10112
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 15838 10112 15844 10124
rect 15620 10084 15665 10112
rect 15799 10084 15844 10112
rect 15620 10072 15626 10084
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 16390 10072 16396 10124
rect 16448 10112 16454 10124
rect 16485 10115 16543 10121
rect 16485 10112 16497 10115
rect 16448 10084 16497 10112
rect 16448 10072 16454 10084
rect 16485 10081 16497 10084
rect 16531 10081 16543 10115
rect 16485 10075 16543 10081
rect 13630 10044 13636 10056
rect 13464 10016 13636 10044
rect 7515 10013 7527 10016
rect 7469 10007 7527 10013
rect 7484 9976 7512 10007
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 7208 9948 7512 9976
rect 8478 9936 8484 9988
rect 8536 9976 8542 9988
rect 9490 9976 9496 9988
rect 8536 9948 9496 9976
rect 8536 9936 8542 9948
rect 9490 9936 9496 9948
rect 9548 9976 9554 9988
rect 10781 9979 10839 9985
rect 10781 9976 10793 9979
rect 9548 9948 10793 9976
rect 9548 9936 9554 9948
rect 10781 9945 10793 9948
rect 10827 9945 10839 9979
rect 10781 9939 10839 9945
rect 12989 9911 13047 9917
rect 12989 9877 13001 9911
rect 13035 9908 13047 9911
rect 13262 9908 13268 9920
rect 13035 9880 13268 9908
rect 13035 9877 13047 9880
rect 12989 9871 13047 9877
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 15286 9908 15292 9920
rect 15247 9880 15292 9908
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 16298 9908 16304 9920
rect 16259 9880 16304 9908
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 1104 9818 17388 9840
rect 1104 9766 3696 9818
rect 3748 9766 3760 9818
rect 3812 9766 3824 9818
rect 3876 9766 3888 9818
rect 3940 9766 9124 9818
rect 9176 9766 9188 9818
rect 9240 9766 9252 9818
rect 9304 9766 9316 9818
rect 9368 9766 14552 9818
rect 14604 9766 14616 9818
rect 14668 9766 14680 9818
rect 14732 9766 14744 9818
rect 14796 9766 17388 9818
rect 1104 9744 17388 9766
rect 5905 9707 5963 9713
rect 5905 9673 5917 9707
rect 5951 9704 5963 9707
rect 15838 9704 15844 9716
rect 5951 9676 6132 9704
rect 5951 9673 5963 9676
rect 5905 9667 5963 9673
rect 6104 9674 6132 9676
rect 7116 9676 7512 9704
rect 15799 9676 15844 9704
rect 6104 9646 6224 9674
rect 5276 9540 5764 9568
rect 5276 9512 5304 9540
rect 3234 9460 3240 9512
rect 3292 9500 3298 9512
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 3292 9472 3617 9500
rect 3292 9460 3298 9472
rect 3605 9469 3617 9472
rect 3651 9500 3663 9503
rect 4617 9503 4675 9509
rect 4617 9500 4629 9503
rect 3651 9472 4629 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 4617 9469 4629 9472
rect 4663 9500 4675 9503
rect 4706 9500 4712 9512
rect 4663 9472 4712 9500
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 5258 9500 5264 9512
rect 5219 9472 5264 9500
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 5736 9509 5764 9540
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9469 5411 9503
rect 5353 9463 5411 9469
rect 5724 9503 5782 9509
rect 5724 9469 5736 9503
rect 5770 9469 5782 9503
rect 5724 9463 5782 9469
rect 5368 9432 5396 9463
rect 6196 9432 6224 9646
rect 6270 9596 6276 9648
rect 6328 9636 6334 9648
rect 7116 9636 7144 9676
rect 6328 9608 7144 9636
rect 6328 9596 6334 9608
rect 7190 9596 7196 9648
rect 7248 9636 7254 9648
rect 7377 9639 7435 9645
rect 7377 9636 7389 9639
rect 7248 9608 7389 9636
rect 7248 9596 7254 9608
rect 7377 9605 7389 9608
rect 7423 9605 7435 9639
rect 7484 9636 7512 9676
rect 15838 9664 15844 9676
rect 15896 9664 15902 9716
rect 7484 9608 7604 9636
rect 7377 9599 7435 9605
rect 7006 9503 7064 9509
rect 7006 9469 7018 9503
rect 7052 9500 7064 9503
rect 7098 9500 7104 9512
rect 7052 9472 7104 9500
rect 7052 9469 7064 9472
rect 7006 9463 7064 9469
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 7466 9500 7472 9512
rect 7427 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7576 9500 7604 9608
rect 10594 9596 10600 9648
rect 10652 9636 10658 9648
rect 10652 9608 11100 9636
rect 10652 9596 10658 9608
rect 9950 9568 9956 9580
rect 9863 9540 9956 9568
rect 9950 9528 9956 9540
rect 10008 9568 10014 9580
rect 11072 9577 11100 9608
rect 12342 9596 12348 9648
rect 12400 9636 12406 9648
rect 12400 9608 13032 9636
rect 12400 9596 12406 9608
rect 13004 9577 13032 9608
rect 10965 9571 11023 9577
rect 10965 9568 10977 9571
rect 10008 9540 10977 9568
rect 10008 9528 10014 9540
rect 8205 9503 8263 9509
rect 8205 9500 8217 9503
rect 7576 9472 8217 9500
rect 8205 9469 8217 9472
rect 8251 9469 8263 9503
rect 10594 9500 10600 9512
rect 10555 9472 10600 9500
rect 8205 9463 8263 9469
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 8481 9435 8539 9441
rect 8481 9432 8493 9435
rect 5368 9404 5764 9432
rect 6196 9404 8493 9432
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3568 9336 3801 9364
rect 3568 9324 3574 9336
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 3789 9327 3847 9333
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 5736 9373 5764 9404
rect 8481 9401 8493 9404
rect 8527 9401 8539 9435
rect 10502 9432 10508 9444
rect 9706 9404 10508 9432
rect 8481 9395 8539 9401
rect 10502 9392 10508 9404
rect 10560 9392 10566 9444
rect 4801 9367 4859 9373
rect 4801 9364 4813 9367
rect 4764 9336 4813 9364
rect 4764 9324 4770 9336
rect 4801 9333 4813 9336
rect 4847 9333 4859 9367
rect 4801 9327 4859 9333
rect 5721 9367 5779 9373
rect 5721 9333 5733 9367
rect 5767 9364 5779 9367
rect 6822 9364 6828 9376
rect 5767 9336 6828 9364
rect 5767 9333 5779 9336
rect 5721 9327 5779 9333
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 7009 9367 7067 9373
rect 7009 9333 7021 9367
rect 7055 9364 7067 9367
rect 7190 9364 7196 9376
rect 7055 9336 7196 9364
rect 7055 9333 7067 9336
rect 7009 9327 7067 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 10410 9364 10416 9376
rect 10371 9336 10416 9364
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 10597 9367 10655 9373
rect 10597 9333 10609 9367
rect 10643 9364 10655 9367
rect 10701 9364 10729 9540
rect 10965 9537 10977 9540
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 13262 9568 13268 9580
rect 13223 9540 13268 9568
rect 12989 9531 13047 9537
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 12434 9500 12440 9512
rect 12299 9472 12440 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 10643 9336 10729 9364
rect 12069 9367 12127 9373
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 12069 9333 12081 9367
rect 12115 9364 12127 9367
rect 12158 9364 12164 9376
rect 12115 9336 12164 9364
rect 12115 9333 12127 9336
rect 12069 9327 12127 9333
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 13004 9364 13032 9531
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9568 14795 9571
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 14783 9540 15301 9568
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 13814 9392 13820 9444
rect 13872 9392 13878 9444
rect 14918 9364 14924 9376
rect 13004 9336 14924 9364
rect 14918 9324 14924 9336
rect 14976 9324 14982 9376
rect 15120 9364 15148 9540
rect 15289 9537 15301 9540
rect 15335 9568 15347 9571
rect 15470 9568 15476 9580
rect 15335 9540 15476 9568
rect 15335 9537 15347 9540
rect 15289 9531 15347 9537
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9500 15255 9503
rect 15562 9500 15568 9512
rect 15243 9472 15568 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 15562 9460 15568 9472
rect 15620 9500 15626 9512
rect 15716 9503 15774 9509
rect 15716 9500 15728 9503
rect 15620 9472 15728 9500
rect 15620 9460 15626 9472
rect 15716 9469 15728 9472
rect 15762 9500 15774 9503
rect 15930 9500 15936 9512
rect 15762 9472 15936 9500
rect 15762 9469 15774 9472
rect 15716 9463 15774 9469
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 15120 9336 15669 9364
rect 15657 9333 15669 9336
rect 15703 9333 15715 9367
rect 15657 9327 15715 9333
rect 1104 9274 17388 9296
rect 1104 9222 6410 9274
rect 6462 9222 6474 9274
rect 6526 9222 6538 9274
rect 6590 9222 6602 9274
rect 6654 9222 11838 9274
rect 11890 9222 11902 9274
rect 11954 9222 11966 9274
rect 12018 9222 12030 9274
rect 12082 9222 17388 9274
rect 1104 9200 17388 9222
rect 1394 9160 1400 9172
rect 1355 9132 1400 9160
rect 1394 9120 1400 9132
rect 1452 9120 1458 9172
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 2682 9160 2688 9172
rect 1627 9132 1992 9160
rect 2643 9132 2688 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 1578 9027 1636 9033
rect 1578 8993 1590 9027
rect 1624 9024 1636 9027
rect 1854 9024 1860 9036
rect 1624 8996 1860 9024
rect 1624 8993 1636 8996
rect 1578 8987 1636 8993
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 1964 8829 1992 9132
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7466 9160 7472 9172
rect 7156 9132 7472 9160
rect 7156 9120 7162 9132
rect 7466 9120 7472 9132
rect 7524 9160 7530 9172
rect 8205 9163 8263 9169
rect 8205 9160 8217 9163
rect 7524 9132 8217 9160
rect 7524 9120 7530 9132
rect 8205 9129 8217 9132
rect 8251 9129 8263 9163
rect 10594 9160 10600 9172
rect 8205 9123 8263 9129
rect 9876 9132 10600 9160
rect 4706 9052 4712 9104
rect 4764 9052 4770 9104
rect 9876 9101 9904 9132
rect 10594 9120 10600 9132
rect 10652 9160 10658 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 10652 9132 12357 9160
rect 10652 9120 10658 9132
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 13170 9160 13176 9172
rect 13131 9132 13176 9160
rect 12345 9123 12403 9129
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 13814 9160 13820 9172
rect 13775 9132 13820 9160
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 15930 9120 15936 9172
rect 15988 9160 15994 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 15988 9132 16681 9160
rect 15988 9120 15994 9132
rect 16669 9129 16681 9132
rect 16715 9129 16727 9163
rect 16669 9123 16727 9129
rect 9861 9095 9919 9101
rect 9861 9061 9873 9095
rect 9907 9061 9919 9095
rect 12158 9092 12164 9104
rect 12098 9064 12164 9092
rect 9861 9055 9919 9061
rect 12158 9052 12164 9064
rect 12216 9052 12222 9104
rect 15197 9095 15255 9101
rect 15197 9061 15209 9095
rect 15243 9092 15255 9095
rect 15286 9092 15292 9104
rect 15243 9064 15292 9092
rect 15243 9061 15255 9064
rect 15197 9055 15255 9061
rect 15286 9052 15292 9064
rect 15344 9052 15350 9104
rect 2590 8984 2596 9036
rect 2648 9024 2654 9036
rect 2682 9027 2740 9033
rect 2682 9024 2694 9027
rect 2648 8996 2694 9024
rect 2648 8984 2654 8996
rect 2682 8993 2694 8996
rect 2728 9024 2740 9027
rect 3145 9027 3203 9033
rect 3145 9024 3157 9027
rect 2728 8996 3157 9024
rect 2728 8993 2740 8996
rect 2682 8987 2740 8993
rect 3145 8993 3157 8996
rect 3191 8993 3203 9027
rect 3145 8987 3203 8993
rect 7834 8984 7840 9036
rect 7892 8984 7898 9036
rect 9585 9027 9643 9033
rect 9585 8993 9597 9027
rect 9631 8993 9643 9027
rect 9766 9024 9772 9036
rect 9727 8996 9772 9024
rect 9585 8987 9643 8993
rect 2038 8916 2044 8968
rect 2096 8956 2102 8968
rect 5721 8959 5779 8965
rect 2096 8928 2141 8956
rect 2096 8916 2102 8928
rect 5721 8925 5733 8959
rect 5767 8956 5779 8959
rect 5997 8959 6055 8965
rect 5767 8928 5948 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8820 2007 8823
rect 2314 8820 2320 8832
rect 1995 8792 2320 8820
rect 1995 8789 2007 8792
rect 1949 8783 2007 8789
rect 2314 8780 2320 8792
rect 2372 8820 2378 8832
rect 2501 8823 2559 8829
rect 2501 8820 2513 8823
rect 2372 8792 2513 8820
rect 2372 8780 2378 8792
rect 2501 8789 2513 8792
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 2682 8780 2688 8832
rect 2740 8820 2746 8832
rect 3053 8823 3111 8829
rect 3053 8820 3065 8823
rect 2740 8792 3065 8820
rect 2740 8780 2746 8792
rect 3053 8789 3065 8792
rect 3099 8820 3111 8823
rect 4249 8823 4307 8829
rect 4249 8820 4261 8823
rect 3099 8792 4261 8820
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 4249 8789 4261 8792
rect 4295 8789 4307 8823
rect 5920 8820 5948 8928
rect 5997 8925 6009 8959
rect 6043 8956 6055 8959
rect 6270 8956 6276 8968
rect 6043 8928 6276 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 6270 8916 6276 8928
rect 6328 8956 6334 8968
rect 6457 8959 6515 8965
rect 6457 8956 6469 8959
rect 6328 8928 6469 8956
rect 6328 8916 6334 8928
rect 6457 8925 6469 8928
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8956 6791 8959
rect 7374 8956 7380 8968
rect 6779 8928 7380 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 9600 8956 9628 8987
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 9950 9024 9956 9036
rect 9911 8996 9956 9024
rect 9950 8984 9956 8996
rect 10008 8984 10014 9036
rect 12986 9024 12992 9036
rect 12947 8996 12992 9024
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13412 8996 13645 9024
rect 13412 8984 13418 8996
rect 13633 8993 13645 8996
rect 13679 8993 13691 9027
rect 14918 9024 14924 9036
rect 14879 8996 14924 9024
rect 13633 8987 13691 8993
rect 14918 8984 14924 8996
rect 14976 8984 14982 9036
rect 16298 8984 16304 9036
rect 16356 8984 16362 9036
rect 10410 8956 10416 8968
rect 9600 8928 10416 8956
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10594 8956 10600 8968
rect 10555 8928 10600 8956
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 10701 8928 10885 8956
rect 10137 8891 10195 8897
rect 10137 8857 10149 8891
rect 10183 8888 10195 8891
rect 10701 8888 10729 8928
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 12802 8956 12808 8968
rect 12715 8928 12808 8956
rect 10873 8919 10931 8925
rect 12802 8916 12808 8928
rect 12860 8956 12866 8968
rect 13722 8956 13728 8968
rect 12860 8928 13728 8956
rect 12860 8916 12866 8928
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 10183 8860 10729 8888
rect 10183 8857 10195 8860
rect 10137 8851 10195 8857
rect 8018 8820 8024 8832
rect 5920 8792 8024 8820
rect 4249 8783 4307 8789
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 1104 8730 17388 8752
rect 1104 8678 3696 8730
rect 3748 8678 3760 8730
rect 3812 8678 3824 8730
rect 3876 8678 3888 8730
rect 3940 8678 9124 8730
rect 9176 8678 9188 8730
rect 9240 8678 9252 8730
rect 9304 8678 9316 8730
rect 9368 8678 14552 8730
rect 14604 8678 14616 8730
rect 14668 8678 14680 8730
rect 14732 8678 14744 8730
rect 14796 8678 17388 8730
rect 1104 8656 17388 8678
rect 2590 8616 2596 8628
rect 2551 8588 2596 8616
rect 2590 8576 2596 8588
rect 2648 8576 2654 8628
rect 6270 8616 6276 8628
rect 4908 8588 6276 8616
rect 4706 8548 4712 8560
rect 4264 8520 4712 8548
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 4264 8480 4292 8520
rect 4706 8508 4712 8520
rect 4764 8508 4770 8560
rect 1903 8452 4292 8480
rect 4341 8483 4399 8489
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4908 8480 4936 8588
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 7374 8616 7380 8628
rect 7335 8588 7380 8616
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 8110 8616 8116 8628
rect 7883 8588 8116 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 9033 8619 9091 8625
rect 9033 8585 9045 8619
rect 9079 8616 9091 8619
rect 9674 8616 9680 8628
rect 9079 8588 9680 8616
rect 9079 8585 9091 8588
rect 9033 8579 9091 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10410 8616 10416 8628
rect 10371 8588 10416 8616
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10560 8588 10977 8616
rect 10560 8576 10566 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12802 8616 12808 8628
rect 12299 8588 12808 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 15105 8619 15163 8625
rect 13280 8588 15056 8616
rect 4985 8551 5043 8557
rect 4985 8517 4997 8551
rect 5031 8548 5043 8551
rect 5442 8548 5448 8560
rect 5031 8520 5448 8548
rect 5031 8517 5043 8520
rect 4985 8511 5043 8517
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 13280 8548 13308 8588
rect 8036 8520 13308 8548
rect 15028 8548 15056 8588
rect 15105 8585 15117 8619
rect 15151 8616 15163 8619
rect 15194 8616 15200 8628
rect 15151 8588 15200 8616
rect 15151 8585 15163 8588
rect 15105 8579 15163 8585
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 15657 8619 15715 8625
rect 15657 8585 15669 8619
rect 15703 8616 15715 8619
rect 15838 8616 15844 8628
rect 15703 8588 15844 8616
rect 15703 8585 15715 8588
rect 15657 8579 15715 8585
rect 15470 8548 15476 8560
rect 15028 8520 15476 8548
rect 7282 8480 7288 8492
rect 4387 8452 4936 8480
rect 5276 8452 7288 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 1670 8412 1676 8424
rect 1631 8384 1676 8412
rect 1670 8372 1676 8384
rect 1728 8372 1734 8424
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 4356 8384 4813 8412
rect 4356 8356 4384 8384
rect 4801 8381 4813 8384
rect 4847 8381 4859 8415
rect 4801 8375 4859 8381
rect 3510 8304 3516 8356
rect 3568 8304 3574 8356
rect 4062 8344 4068 8356
rect 4023 8316 4068 8344
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 4338 8304 4344 8356
rect 4396 8304 4402 8356
rect 4706 8304 4712 8356
rect 4764 8344 4770 8356
rect 5276 8344 5304 8452
rect 7282 8440 7288 8452
rect 7340 8480 7346 8492
rect 7340 8452 7420 8480
rect 7340 8440 7346 8452
rect 5442 8372 5448 8424
rect 5500 8412 5506 8424
rect 5629 8415 5687 8421
rect 5629 8412 5641 8415
rect 5500 8384 5641 8412
rect 5500 8372 5506 8384
rect 5629 8381 5641 8384
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 5810 8372 5816 8424
rect 5868 8412 5874 8424
rect 6089 8415 6147 8421
rect 6089 8412 6101 8415
rect 5868 8384 6101 8412
rect 5868 8372 5874 8384
rect 6089 8381 6101 8384
rect 6135 8381 6147 8415
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 6089 8375 6147 8381
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 7098 8412 7104 8424
rect 7059 8384 7104 8412
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 7248 8384 7293 8412
rect 7248 8372 7254 8384
rect 4764 8316 5304 8344
rect 4764 8304 4770 8316
rect 1489 8279 1547 8285
rect 1489 8245 1501 8279
rect 1535 8276 1547 8279
rect 2038 8276 2044 8288
rect 1535 8248 2044 8276
rect 1535 8245 1547 8248
rect 1489 8239 1547 8245
rect 2038 8236 2044 8248
rect 2096 8276 2102 8288
rect 2498 8276 2504 8288
rect 2096 8248 2504 8276
rect 2096 8236 2102 8248
rect 2498 8236 2504 8248
rect 2556 8236 2562 8288
rect 5276 8276 5304 8316
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 7009 8347 7067 8353
rect 7009 8344 7021 8347
rect 5408 8316 7021 8344
rect 5408 8304 5414 8316
rect 7009 8313 7021 8316
rect 7055 8313 7067 8347
rect 7392 8344 7420 8452
rect 8036 8421 8064 8520
rect 15470 8508 15476 8520
rect 15528 8508 15534 8560
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 8812 8452 11192 8480
rect 8812 8440 8818 8452
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 8113 8415 8171 8421
rect 8113 8381 8125 8415
rect 8159 8412 8171 8415
rect 8665 8415 8723 8421
rect 8665 8412 8677 8415
rect 8159 8384 8677 8412
rect 8159 8381 8171 8384
rect 8113 8375 8171 8381
rect 8665 8381 8677 8384
rect 8711 8381 8723 8415
rect 8665 8375 8723 8381
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8381 8907 8415
rect 8849 8375 8907 8381
rect 8128 8344 8156 8375
rect 7392 8316 8156 8344
rect 7009 8307 7067 8313
rect 8570 8304 8576 8356
rect 8628 8344 8634 8356
rect 8864 8344 8892 8375
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 10014 8415 10072 8421
rect 10014 8412 10026 8415
rect 9824 8384 10026 8412
rect 9824 8372 9830 8384
rect 10014 8381 10026 8384
rect 10060 8412 10072 8415
rect 10502 8412 10508 8424
rect 10060 8384 10508 8412
rect 10060 8381 10072 8384
rect 10014 8375 10072 8381
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 11164 8421 11192 8452
rect 13538 8440 13544 8492
rect 13596 8480 13602 8492
rect 14277 8483 14335 8489
rect 14277 8480 14289 8483
rect 13596 8452 14289 8480
rect 13596 8440 13602 8452
rect 14277 8449 14289 8452
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8480 14611 8483
rect 14918 8480 14924 8492
rect 14599 8452 14924 8480
rect 14599 8449 14611 8452
rect 14553 8443 14611 8449
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 12069 8415 12127 8421
rect 12069 8381 12081 8415
rect 12115 8412 12127 8415
rect 12158 8412 12164 8424
rect 12115 8384 12164 8412
rect 12115 8381 12127 8384
rect 12069 8375 12127 8381
rect 12158 8372 12164 8384
rect 12216 8372 12222 8424
rect 15258 8415 15316 8421
rect 15258 8381 15270 8415
rect 15304 8412 15316 8415
rect 15562 8412 15568 8424
rect 15304 8384 15568 8412
rect 15304 8381 15316 8384
rect 15258 8375 15316 8381
rect 15562 8372 15568 8384
rect 15620 8372 15626 8424
rect 8628 8316 8892 8344
rect 10110 8347 10168 8353
rect 8628 8304 8634 8316
rect 10110 8313 10122 8347
rect 10156 8344 10168 8347
rect 10410 8344 10416 8356
rect 10156 8316 10416 8344
rect 10156 8313 10168 8316
rect 10110 8307 10168 8313
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 13814 8304 13820 8356
rect 13872 8304 13878 8356
rect 15354 8347 15412 8353
rect 15354 8313 15366 8347
rect 15400 8344 15412 8347
rect 15672 8344 15700 8579
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 15746 8508 15752 8560
rect 15804 8508 15810 8560
rect 15764 8421 15792 8508
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8381 15807 8415
rect 16390 8412 16396 8424
rect 16351 8384 16396 8412
rect 15749 8375 15807 8381
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 15400 8316 15700 8344
rect 15400 8313 15412 8316
rect 15354 8307 15412 8313
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5276 8248 5457 8276
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 6270 8276 6276 8288
rect 6183 8248 6276 8276
rect 5445 8239 5503 8245
rect 6270 8236 6276 8248
rect 6328 8276 6334 8288
rect 6730 8276 6736 8288
rect 6328 8248 6736 8276
rect 6328 8236 6334 8248
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 9861 8279 9919 8285
rect 9861 8245 9873 8279
rect 9907 8276 9919 8279
rect 9950 8276 9956 8288
rect 9907 8248 9956 8276
rect 9907 8245 9919 8248
rect 9861 8239 9919 8245
rect 9950 8236 9956 8248
rect 10008 8236 10014 8288
rect 10594 8236 10600 8288
rect 10652 8276 10658 8288
rect 12342 8276 12348 8288
rect 10652 8248 12348 8276
rect 10652 8236 10658 8248
rect 12342 8236 12348 8248
rect 12400 8236 12406 8288
rect 12802 8276 12808 8288
rect 12763 8248 12808 8276
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 15838 8236 15844 8288
rect 15896 8276 15902 8288
rect 16209 8279 16267 8285
rect 16209 8276 16221 8279
rect 15896 8248 16221 8276
rect 15896 8236 15902 8248
rect 16209 8245 16221 8248
rect 16255 8245 16267 8279
rect 16209 8239 16267 8245
rect 1104 8186 17388 8208
rect 1104 8134 6410 8186
rect 6462 8134 6474 8186
rect 6526 8134 6538 8186
rect 6590 8134 6602 8186
rect 6654 8134 11838 8186
rect 11890 8134 11902 8186
rect 11954 8134 11966 8186
rect 12018 8134 12030 8186
rect 12082 8134 17388 8186
rect 1104 8112 17388 8134
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 1765 8075 1823 8081
rect 1765 8072 1777 8075
rect 1728 8044 1777 8072
rect 1728 8032 1734 8044
rect 1765 8041 1777 8044
rect 1811 8041 1823 8075
rect 1765 8035 1823 8041
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 4062 8072 4068 8084
rect 2915 8044 4068 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 5408 8044 5457 8072
rect 5408 8032 5414 8044
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 11054 8072 11060 8084
rect 5445 8035 5503 8041
rect 8036 8044 11060 8072
rect 2590 8004 2596 8016
rect 2551 7976 2596 8004
rect 2590 7964 2596 7976
rect 2648 7964 2654 8016
rect 4614 8004 4620 8016
rect 4448 7976 4620 8004
rect 1946 7936 1952 7948
rect 1907 7908 1952 7936
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 2314 7936 2320 7948
rect 2275 7908 2320 7936
rect 2314 7896 2320 7908
rect 2372 7896 2378 7948
rect 2498 7936 2504 7948
rect 2459 7908 2504 7936
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 2682 7936 2688 7948
rect 2643 7908 2688 7936
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 4448 7945 4476 7976
rect 4614 7964 4620 7976
rect 4672 7964 4678 8016
rect 7834 7964 7840 8016
rect 7892 8004 7898 8016
rect 8036 8013 8064 8044
rect 11054 8032 11060 8044
rect 11112 8072 11118 8084
rect 11517 8075 11575 8081
rect 11112 8044 11376 8072
rect 11112 8032 11118 8044
rect 8021 8007 8079 8013
rect 8021 8004 8033 8007
rect 7892 7976 8033 8004
rect 7892 7964 7898 7976
rect 8021 7973 8033 7976
rect 8067 7973 8079 8007
rect 8021 7967 8079 7973
rect 8205 8007 8263 8013
rect 8205 7973 8217 8007
rect 8251 8004 8263 8007
rect 8754 8004 8760 8016
rect 8251 7976 8760 8004
rect 8251 7973 8263 7976
rect 8205 7967 8263 7973
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 9950 7964 9956 8016
rect 10008 8004 10014 8016
rect 10045 8007 10103 8013
rect 10045 8004 10057 8007
rect 10008 7976 10057 8004
rect 10008 7964 10014 7976
rect 10045 7973 10057 7976
rect 10091 7973 10103 8007
rect 10045 7967 10103 7973
rect 10778 7964 10784 8016
rect 10836 7964 10842 8016
rect 11348 8004 11376 8044
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 12161 8075 12219 8081
rect 12161 8072 12173 8075
rect 11563 8044 12173 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 12161 8041 12173 8044
rect 12207 8072 12219 8075
rect 12526 8072 12532 8084
rect 12207 8044 12532 8072
rect 12207 8041 12219 8044
rect 12161 8035 12219 8041
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 13814 8072 13820 8084
rect 13775 8044 13820 8072
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 14918 8072 14924 8084
rect 14879 8044 14924 8072
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 15565 8075 15623 8081
rect 15565 8041 15577 8075
rect 15611 8072 15623 8075
rect 15654 8072 15660 8084
rect 15611 8044 15660 8072
rect 15611 8041 15623 8044
rect 15565 8035 15623 8041
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 12434 8004 12440 8016
rect 11348 7976 12440 8004
rect 12434 7964 12440 7976
rect 12492 8004 12498 8016
rect 13170 8004 13176 8016
rect 12492 7976 13176 8004
rect 12492 7964 12498 7976
rect 13170 7964 13176 7976
rect 13228 8004 13234 8016
rect 13228 7976 13676 8004
rect 13228 7964 13234 7976
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7905 4491 7939
rect 4433 7899 4491 7905
rect 4522 7896 4528 7948
rect 4580 7936 4586 7948
rect 4580 7908 4625 7936
rect 4580 7896 4586 7908
rect 4706 7896 4712 7948
rect 4764 7936 4770 7948
rect 5261 7939 5319 7945
rect 5261 7936 5273 7939
rect 4764 7908 5273 7936
rect 4764 7896 4770 7908
rect 5261 7905 5273 7908
rect 5307 7905 5319 7939
rect 9490 7936 9496 7948
rect 9451 7908 9496 7936
rect 5261 7899 5319 7905
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 13648 7945 13676 7976
rect 13722 7964 13728 8016
rect 13780 8004 13786 8016
rect 13780 7976 15884 8004
rect 13780 7964 13786 7976
rect 12158 7939 12216 7945
rect 12158 7905 12170 7939
rect 12204 7936 12216 7939
rect 13633 7939 13691 7945
rect 12204 7908 12434 7936
rect 12204 7905 12216 7908
rect 12158 7899 12216 7905
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5442 7868 5448 7880
rect 5123 7840 5448 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7868 9827 7871
rect 10594 7868 10600 7880
rect 9815 7840 10600 7868
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 12406 7868 12434 7908
rect 13633 7905 13645 7939
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 14737 7939 14795 7945
rect 14737 7905 14749 7939
rect 14783 7905 14795 7939
rect 14737 7899 14795 7905
rect 12621 7871 12679 7877
rect 12621 7868 12633 7871
rect 12406 7840 12633 7868
rect 12621 7837 12633 7840
rect 12667 7868 12679 7871
rect 12802 7868 12808 7880
rect 12667 7840 12808 7868
rect 12667 7837 12679 7840
rect 12621 7831 12679 7837
rect 12802 7828 12808 7840
rect 12860 7868 12866 7880
rect 13078 7868 13084 7880
rect 12860 7840 13084 7868
rect 12860 7828 12866 7840
rect 13078 7828 13084 7840
rect 13136 7828 13142 7880
rect 12250 7760 12256 7812
rect 12308 7800 12314 7812
rect 14752 7800 14780 7899
rect 15286 7896 15292 7948
rect 15344 7936 15350 7948
rect 15856 7945 15884 7976
rect 15749 7939 15807 7945
rect 15749 7936 15761 7939
rect 15344 7908 15761 7936
rect 15344 7896 15350 7908
rect 15749 7905 15761 7908
rect 15795 7905 15807 7939
rect 15749 7899 15807 7905
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7905 15899 7939
rect 16666 7936 16672 7948
rect 16627 7908 16672 7936
rect 15841 7899 15899 7905
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 12308 7772 14780 7800
rect 12308 7760 12314 7772
rect 15470 7760 15476 7812
rect 15528 7800 15534 7812
rect 16485 7803 16543 7809
rect 16485 7800 16497 7803
rect 15528 7772 16497 7800
rect 15528 7760 15534 7772
rect 16485 7769 16497 7772
rect 16531 7769 16543 7803
rect 16485 7763 16543 7769
rect 4246 7732 4252 7744
rect 4207 7704 4252 7732
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 9674 7732 9680 7744
rect 9587 7704 9680 7732
rect 9674 7692 9680 7704
rect 9732 7732 9738 7744
rect 10410 7732 10416 7744
rect 9732 7704 10416 7732
rect 9732 7692 9738 7704
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 11977 7735 12035 7741
rect 11977 7701 11989 7735
rect 12023 7732 12035 7735
rect 12158 7732 12164 7744
rect 12023 7704 12164 7732
rect 12023 7701 12035 7704
rect 11977 7695 12035 7701
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 12526 7732 12532 7744
rect 12439 7704 12532 7732
rect 12526 7692 12532 7704
rect 12584 7732 12590 7744
rect 13354 7732 13360 7744
rect 12584 7704 13360 7732
rect 12584 7692 12590 7704
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 1104 7642 17388 7664
rect 1104 7590 3696 7642
rect 3748 7590 3760 7642
rect 3812 7590 3824 7642
rect 3876 7590 3888 7642
rect 3940 7590 9124 7642
rect 9176 7590 9188 7642
rect 9240 7590 9252 7642
rect 9304 7590 9316 7642
rect 9368 7590 14552 7642
rect 14604 7590 14616 7642
rect 14668 7590 14680 7642
rect 14732 7590 14744 7642
rect 14796 7590 17388 7642
rect 1104 7568 17388 7590
rect 2593 7531 2651 7537
rect 2593 7497 2605 7531
rect 2639 7528 2651 7531
rect 2639 7500 3188 7528
rect 2639 7497 2651 7500
rect 2593 7491 2651 7497
rect 2608 7460 2636 7491
rect 3160 7469 3188 7500
rect 3510 7488 3516 7540
rect 3568 7528 3574 7540
rect 3697 7531 3755 7537
rect 3697 7528 3709 7531
rect 3568 7500 3709 7528
rect 3568 7488 3574 7500
rect 3697 7497 3709 7500
rect 3743 7528 3755 7531
rect 4062 7528 4068 7540
rect 3743 7500 4068 7528
rect 3743 7497 3755 7500
rect 3697 7491 3755 7497
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 10502 7528 10508 7540
rect 5500 7500 9812 7528
rect 10463 7500 10508 7528
rect 5500 7488 5506 7500
rect 3145 7463 3203 7469
rect 2148 7432 2636 7460
rect 2700 7432 3096 7460
rect 1670 7148 1676 7200
rect 1728 7188 1734 7200
rect 2041 7191 2099 7197
rect 2041 7188 2053 7191
rect 1728 7160 2053 7188
rect 1728 7148 1734 7160
rect 2041 7157 2053 7160
rect 2087 7157 2099 7191
rect 2148 7188 2176 7432
rect 2700 7401 2728 7432
rect 2685 7395 2743 7401
rect 2685 7392 2697 7395
rect 2516 7364 2697 7392
rect 2222 7327 2280 7333
rect 2222 7293 2234 7327
rect 2268 7324 2280 7327
rect 2516 7324 2544 7364
rect 2685 7361 2697 7364
rect 2731 7361 2743 7395
rect 3068 7392 3096 7432
rect 3145 7429 3157 7463
rect 3191 7460 3203 7463
rect 3191 7432 4844 7460
rect 3191 7429 3203 7432
rect 3145 7423 3203 7429
rect 4246 7392 4252 7404
rect 3068 7364 4252 7392
rect 2685 7355 2743 7361
rect 4246 7352 4252 7364
rect 4304 7392 4310 7404
rect 4304 7364 4660 7392
rect 4304 7352 4310 7364
rect 2268 7296 2544 7324
rect 2268 7293 2280 7296
rect 2222 7287 2280 7293
rect 3142 7284 3148 7336
rect 3200 7324 3206 7336
rect 3270 7327 3328 7333
rect 3270 7324 3282 7327
rect 3200 7296 3282 7324
rect 3200 7284 3206 7296
rect 3270 7293 3282 7296
rect 3316 7324 3328 7327
rect 3789 7327 3847 7333
rect 3316 7296 3648 7324
rect 3316 7293 3328 7296
rect 3270 7287 3328 7293
rect 3620 7256 3648 7296
rect 3789 7293 3801 7327
rect 3835 7293 3847 7327
rect 3789 7287 3847 7293
rect 3804 7256 3832 7287
rect 4062 7284 4068 7336
rect 4120 7324 4126 7336
rect 4632 7333 4660 7364
rect 4816 7333 4844 7432
rect 5810 7420 5816 7472
rect 5868 7460 5874 7472
rect 7469 7463 7527 7469
rect 7469 7460 7481 7463
rect 5868 7432 7481 7460
rect 5868 7420 5874 7432
rect 7469 7429 7481 7432
rect 7515 7429 7527 7463
rect 7469 7423 7527 7429
rect 7650 7420 7656 7472
rect 7708 7460 7714 7472
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 7708 7432 7849 7460
rect 7708 7420 7714 7432
rect 7837 7429 7849 7432
rect 7883 7429 7895 7463
rect 7837 7423 7895 7429
rect 8478 7420 8484 7472
rect 8536 7460 8542 7472
rect 8941 7463 8999 7469
rect 8941 7460 8953 7463
rect 8536 7432 8953 7460
rect 8536 7420 8542 7432
rect 8941 7429 8953 7432
rect 8987 7429 8999 7463
rect 8941 7423 8999 7429
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 5905 7395 5963 7401
rect 5905 7392 5917 7395
rect 5776 7364 5917 7392
rect 5776 7352 5782 7364
rect 5905 7361 5917 7364
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 9674 7392 9680 7404
rect 7791 7364 8248 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 4433 7327 4491 7333
rect 4433 7324 4445 7327
rect 4120 7296 4445 7324
rect 4120 7284 4126 7296
rect 4433 7293 4445 7296
rect 4479 7293 4491 7327
rect 4433 7287 4491 7293
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 5442 7327 5500 7333
rect 5442 7293 5454 7327
rect 5488 7324 5500 7327
rect 5736 7324 5764 7352
rect 8220 7336 8248 7364
rect 8309 7364 9680 7392
rect 5488 7296 5764 7324
rect 5813 7327 5871 7333
rect 5488 7293 5500 7296
rect 5442 7287 5500 7293
rect 5813 7293 5825 7327
rect 5859 7293 5871 7327
rect 7006 7324 7012 7336
rect 6967 7296 7012 7324
rect 5813 7287 5871 7293
rect 4525 7259 4583 7265
rect 4525 7256 4537 7259
rect 3620 7228 4537 7256
rect 4525 7225 4537 7228
rect 4571 7225 4583 7259
rect 5828 7256 5856 7287
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7293 7711 7327
rect 8202 7324 8208 7336
rect 8115 7296 8208 7324
rect 7653 7287 7711 7293
rect 4525 7219 4583 7225
rect 5460 7228 5856 7256
rect 7668 7256 7696 7287
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8309 7256 8337 7364
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 9784 7392 9812 7500
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 10778 7488 10784 7540
rect 10836 7528 10842 7540
rect 10965 7531 11023 7537
rect 10965 7528 10977 7531
rect 10836 7500 10977 7528
rect 10836 7488 10842 7500
rect 10965 7497 10977 7500
rect 11011 7497 11023 7531
rect 15657 7531 15715 7537
rect 15657 7528 15669 7531
rect 10965 7491 11023 7497
rect 12406 7500 15669 7528
rect 12406 7460 12434 7500
rect 15657 7497 15669 7500
rect 15703 7497 15715 7531
rect 15657 7491 15715 7497
rect 12176 7432 12434 7460
rect 10137 7395 10195 7401
rect 10137 7392 10149 7395
rect 9784 7364 10149 7392
rect 10137 7361 10149 7364
rect 10183 7392 10195 7395
rect 12066 7392 12072 7404
rect 10183 7364 12072 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 8846 7324 8852 7336
rect 8759 7296 8852 7324
rect 8846 7284 8852 7296
rect 8904 7324 8910 7336
rect 9368 7327 9426 7333
rect 9368 7324 9380 7327
rect 8904 7296 9380 7324
rect 8904 7284 8910 7296
rect 9368 7293 9380 7296
rect 9414 7324 9426 7327
rect 10318 7324 10324 7336
rect 9414 7296 9720 7324
rect 10279 7296 10324 7324
rect 9414 7293 9426 7296
rect 9368 7287 9426 7293
rect 7668 7228 8337 7256
rect 9692 7256 9720 7296
rect 10318 7284 10324 7296
rect 10376 7284 10382 7336
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 11112 7296 11161 7324
rect 11112 7284 11118 7296
rect 11149 7293 11161 7296
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 12176 7256 12204 7432
rect 16206 7392 16212 7404
rect 12268 7364 16212 7392
rect 12268 7333 12296 7364
rect 16206 7352 16212 7364
rect 16264 7352 16270 7404
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7293 12311 7327
rect 12253 7287 12311 7293
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 12989 7327 13047 7333
rect 12989 7324 13001 7327
rect 12400 7296 13001 7324
rect 12400 7284 12406 7296
rect 12989 7293 13001 7296
rect 13035 7293 13047 7327
rect 15838 7324 15844 7336
rect 15799 7296 15844 7324
rect 12989 7287 13047 7293
rect 15838 7284 15844 7296
rect 15896 7284 15902 7336
rect 15930 7284 15936 7336
rect 15988 7324 15994 7336
rect 15988 7296 16033 7324
rect 15988 7284 15994 7296
rect 13262 7256 13268 7268
rect 9692 7228 12204 7256
rect 13223 7228 13268 7256
rect 5460 7200 5488 7228
rect 13262 7216 13268 7228
rect 13320 7216 13326 7268
rect 13814 7216 13820 7268
rect 13872 7216 13878 7268
rect 2225 7191 2283 7197
rect 2225 7188 2237 7191
rect 2148 7160 2237 7188
rect 2041 7151 2099 7157
rect 2225 7157 2237 7160
rect 2271 7157 2283 7191
rect 2225 7151 2283 7157
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7188 3387 7191
rect 3510 7188 3516 7200
rect 3375 7160 3516 7188
rect 3375 7157 3387 7160
rect 3329 7151 3387 7157
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 4246 7188 4252 7200
rect 4207 7160 4252 7188
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 4798 7148 4804 7200
rect 4856 7188 4862 7200
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 4856 7160 5273 7188
rect 4856 7148 4862 7160
rect 5261 7157 5273 7160
rect 5307 7157 5319 7191
rect 5442 7188 5448 7200
rect 5403 7160 5448 7188
rect 5261 7151 5319 7157
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6144 7160 6837 7188
rect 6144 7148 6150 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 6825 7151 6883 7157
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 8205 7191 8263 7197
rect 8205 7188 8217 7191
rect 7708 7160 8217 7188
rect 7708 7148 7714 7160
rect 8205 7157 8217 7160
rect 8251 7157 8263 7191
rect 8205 7151 8263 7157
rect 8389 7191 8447 7197
rect 8389 7157 8401 7191
rect 8435 7188 8447 7191
rect 8478 7188 8484 7200
rect 8435 7160 8484 7188
rect 8435 7157 8447 7160
rect 8389 7151 8447 7157
rect 8478 7148 8484 7160
rect 8536 7188 8542 7200
rect 9309 7191 9367 7197
rect 9309 7188 9321 7191
rect 8536 7160 9321 7188
rect 8536 7148 8542 7160
rect 9309 7157 9321 7160
rect 9355 7157 9367 7191
rect 9490 7188 9496 7200
rect 9451 7160 9496 7188
rect 9309 7151 9367 7157
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 14737 7191 14795 7197
rect 12492 7160 12537 7188
rect 12492 7148 12498 7160
rect 14737 7157 14749 7191
rect 14783 7188 14795 7191
rect 15010 7188 15016 7200
rect 14783 7160 15016 7188
rect 14783 7157 14795 7160
rect 14737 7151 14795 7157
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 1104 7098 17388 7120
rect 1104 7046 6410 7098
rect 6462 7046 6474 7098
rect 6526 7046 6538 7098
rect 6590 7046 6602 7098
rect 6654 7046 11838 7098
rect 11890 7046 11902 7098
rect 11954 7046 11966 7098
rect 12018 7046 12030 7098
rect 12082 7046 17388 7098
rect 1104 7024 17388 7046
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7064 6956 8892 6984
rect 7064 6944 7070 6956
rect 1670 6916 1676 6928
rect 1631 6888 1676 6916
rect 1670 6876 1676 6888
rect 1728 6876 1734 6928
rect 2406 6876 2412 6928
rect 2464 6876 2470 6928
rect 4798 6916 4804 6928
rect 4759 6888 4804 6916
rect 4798 6876 4804 6888
rect 4856 6876 4862 6928
rect 6086 6916 6092 6928
rect 6026 6888 6092 6916
rect 6086 6876 6092 6888
rect 6144 6876 6150 6928
rect 8234 6888 8800 6916
rect 6730 6848 6736 6860
rect 6691 6820 6736 6848
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6780 1455 6783
rect 2038 6780 2044 6792
rect 1443 6752 2044 6780
rect 1443 6749 1455 6752
rect 1397 6743 1455 6749
rect 2038 6740 2044 6752
rect 2096 6740 2102 6792
rect 2314 6740 2320 6792
rect 2372 6780 2378 6792
rect 3145 6783 3203 6789
rect 3145 6780 3157 6783
rect 2372 6752 3157 6780
rect 2372 6740 2378 6752
rect 3145 6749 3157 6752
rect 3191 6749 3203 6783
rect 3145 6743 3203 6749
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 4890 6780 4896 6792
rect 4571 6752 4896 6780
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 7006 6780 7012 6792
rect 6967 6752 7012 6780
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 8260 6752 8493 6780
rect 8260 6740 8266 6752
rect 8481 6749 8493 6752
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 8772 6712 8800 6888
rect 8864 6848 8892 6956
rect 12158 6944 12164 6996
rect 12216 6984 12222 6996
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 12216 6956 12357 6984
rect 12216 6944 12222 6956
rect 12345 6953 12357 6956
rect 12391 6953 12403 6987
rect 12345 6947 12403 6953
rect 12529 6987 12587 6993
rect 12529 6953 12541 6987
rect 12575 6984 12587 6987
rect 13262 6984 13268 6996
rect 12575 6956 13268 6984
rect 12575 6953 12587 6956
rect 12529 6947 12587 6953
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 13173 6919 13231 6925
rect 13173 6916 13185 6919
rect 12452 6888 13185 6916
rect 12452 6860 12480 6888
rect 13173 6885 13185 6888
rect 13219 6885 13231 6919
rect 13173 6879 13231 6885
rect 9493 6851 9551 6857
rect 9493 6848 9505 6851
rect 8864 6820 9505 6848
rect 9493 6817 9505 6820
rect 9539 6848 9551 6851
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 9539 6820 10333 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 10321 6811 10379 6817
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 10781 6851 10839 6857
rect 10781 6848 10793 6851
rect 10468 6820 10793 6848
rect 10468 6808 10474 6820
rect 10781 6817 10793 6820
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 11885 6851 11943 6857
rect 11885 6817 11897 6851
rect 11931 6848 11943 6851
rect 12348 6851 12406 6857
rect 12348 6848 12360 6851
rect 11931 6820 12360 6848
rect 11931 6817 11943 6820
rect 11885 6811 11943 6817
rect 12348 6817 12360 6820
rect 12394 6848 12406 6851
rect 12434 6848 12440 6860
rect 12394 6820 12440 6848
rect 12394 6817 12406 6820
rect 12348 6811 12406 6817
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12158 6780 12164 6792
rect 12023 6752 12164 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12158 6740 12164 6752
rect 12216 6780 12222 6792
rect 13004 6780 13032 6811
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 13136 6820 13277 6848
rect 13136 6808 13142 6820
rect 13265 6817 13277 6820
rect 13311 6817 13323 6851
rect 13265 6811 13323 6817
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 13412 6820 13457 6848
rect 13412 6808 13418 6820
rect 14918 6808 14924 6860
rect 14976 6848 14982 6860
rect 15105 6851 15163 6857
rect 15105 6848 15117 6851
rect 14976 6820 15117 6848
rect 14976 6808 14982 6820
rect 15105 6817 15117 6820
rect 15151 6817 15163 6851
rect 15105 6811 15163 6817
rect 15289 6851 15347 6857
rect 15289 6817 15301 6851
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 12216 6752 13032 6780
rect 12216 6740 12222 6752
rect 10137 6715 10195 6721
rect 10137 6712 10149 6715
rect 8772 6684 10149 6712
rect 10137 6681 10149 6684
rect 10183 6681 10195 6715
rect 10137 6675 10195 6681
rect 10594 6672 10600 6724
rect 10652 6712 10658 6724
rect 13538 6712 13544 6724
rect 10652 6684 13400 6712
rect 13499 6684 13544 6712
rect 10652 6672 10658 6684
rect 6273 6647 6331 6653
rect 6273 6613 6285 6647
rect 6319 6644 6331 6647
rect 7650 6644 7656 6656
rect 6319 6616 7656 6644
rect 6319 6613 6331 6616
rect 6273 6607 6331 6613
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 9677 6647 9735 6653
rect 9677 6613 9689 6647
rect 9723 6644 9735 6647
rect 9766 6644 9772 6656
rect 9723 6616 9772 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 10965 6647 11023 6653
rect 10965 6613 10977 6647
rect 11011 6644 11023 6647
rect 12250 6644 12256 6656
rect 11011 6616 12256 6644
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 13372 6644 13400 6684
rect 13538 6672 13544 6684
rect 13596 6672 13602 6724
rect 14366 6672 14372 6724
rect 14424 6712 14430 6724
rect 15304 6712 15332 6811
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 15562 6857 15568 6860
rect 15519 6851 15568 6857
rect 15436 6820 15481 6848
rect 15436 6808 15442 6820
rect 15519 6817 15531 6851
rect 15565 6817 15568 6851
rect 15519 6811 15568 6817
rect 15562 6808 15568 6811
rect 15620 6808 15626 6860
rect 16114 6808 16120 6860
rect 16172 6848 16178 6860
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 16172 6820 16313 6848
rect 16172 6808 16178 6820
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 16301 6811 16359 6817
rect 15654 6740 15660 6792
rect 15712 6780 15718 6792
rect 15930 6780 15936 6792
rect 15712 6752 15936 6780
rect 15712 6740 15718 6752
rect 15930 6740 15936 6752
rect 15988 6780 15994 6792
rect 16485 6783 16543 6789
rect 16485 6780 16497 6783
rect 15988 6752 16497 6780
rect 15988 6740 15994 6752
rect 16485 6749 16497 6752
rect 16531 6749 16543 6783
rect 16485 6743 16543 6749
rect 16117 6715 16175 6721
rect 16117 6712 16129 6715
rect 14424 6684 16129 6712
rect 14424 6672 14430 6684
rect 16117 6681 16129 6684
rect 16163 6681 16175 6715
rect 16117 6675 16175 6681
rect 15102 6644 15108 6656
rect 13372 6616 15108 6644
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 15194 6604 15200 6656
rect 15252 6644 15258 6656
rect 15657 6647 15715 6653
rect 15657 6644 15669 6647
rect 15252 6616 15669 6644
rect 15252 6604 15258 6616
rect 15657 6613 15669 6616
rect 15703 6613 15715 6647
rect 15657 6607 15715 6613
rect 1104 6554 17388 6576
rect 1104 6502 3696 6554
rect 3748 6502 3760 6554
rect 3812 6502 3824 6554
rect 3876 6502 3888 6554
rect 3940 6502 9124 6554
rect 9176 6502 9188 6554
rect 9240 6502 9252 6554
rect 9304 6502 9316 6554
rect 9368 6502 14552 6554
rect 14604 6502 14616 6554
rect 14668 6502 14680 6554
rect 14732 6502 14744 6554
rect 14796 6502 17388 6554
rect 1104 6480 17388 6502
rect 2406 6440 2412 6452
rect 2367 6412 2412 6440
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 3142 6440 3148 6452
rect 3103 6412 3148 6440
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 7006 6400 7012 6452
rect 7064 6440 7070 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7064 6412 7941 6440
rect 7064 6400 7070 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 11146 6440 11152 6452
rect 7929 6403 7987 6409
rect 8036 6412 11152 6440
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 4617 6307 4675 6313
rect 4617 6304 4629 6307
rect 4304 6276 4629 6304
rect 4304 6264 4310 6276
rect 4617 6273 4629 6276
rect 4663 6273 4675 6307
rect 8036 6304 8064 6412
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 13814 6440 13820 6452
rect 13403 6412 13820 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 13909 6443 13967 6449
rect 13909 6409 13921 6443
rect 13955 6440 13967 6443
rect 14918 6440 14924 6452
rect 13955 6412 14924 6440
rect 13955 6409 13967 6412
rect 13909 6403 13967 6409
rect 4617 6267 4675 6273
rect 5460 6276 8064 6304
rect 9309 6307 9367 6313
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2774 6236 2780 6248
rect 2271 6208 2780 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 4890 6196 4896 6248
rect 4948 6236 4954 6248
rect 4948 6208 4993 6236
rect 4948 6196 4954 6208
rect 5166 6196 5172 6248
rect 5224 6236 5230 6248
rect 5353 6239 5411 6245
rect 5353 6236 5365 6239
rect 5224 6208 5365 6236
rect 5224 6196 5230 6208
rect 5353 6205 5365 6208
rect 5399 6205 5411 6239
rect 5353 6199 5411 6205
rect 4154 6128 4160 6180
rect 4212 6128 4218 6180
rect 1578 6060 1584 6112
rect 1636 6100 1642 6112
rect 5460 6100 5488 6276
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9398 6304 9404 6316
rect 9355 6276 9404 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 5537 6239 5595 6245
rect 5537 6205 5549 6239
rect 5583 6236 5595 6239
rect 5626 6236 5632 6248
rect 5583 6208 5632 6236
rect 5583 6205 5595 6208
rect 5537 6199 5595 6205
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 7098 6236 7104 6248
rect 7059 6208 7104 6236
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7708 6208 8125 6236
rect 7708 6196 7714 6208
rect 8113 6205 8125 6208
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 8202 6196 8208 6248
rect 8260 6236 8266 6248
rect 8478 6236 8484 6248
rect 8260 6208 8305 6236
rect 8439 6208 8484 6236
rect 8260 6196 8266 6208
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6205 9091 6239
rect 9033 6199 9091 6205
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6236 12127 6239
rect 12250 6236 12256 6248
rect 12115 6208 12256 6236
rect 12115 6205 12127 6208
rect 12069 6199 12127 6205
rect 8297 6171 8355 6177
rect 8297 6137 8309 6171
rect 8343 6168 8355 6171
rect 8846 6168 8852 6180
rect 8343 6140 8852 6168
rect 8343 6137 8355 6140
rect 8297 6131 8355 6137
rect 8846 6128 8852 6140
rect 8904 6128 8910 6180
rect 5718 6100 5724 6112
rect 1636 6072 5488 6100
rect 5679 6072 5724 6100
rect 1636 6060 1642 6072
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 6914 6100 6920 6112
rect 6875 6072 6920 6100
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 9048 6100 9076 6199
rect 12250 6196 12256 6208
rect 12308 6196 12314 6248
rect 13170 6236 13176 6248
rect 13131 6208 13176 6236
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 14366 6245 14372 6248
rect 13817 6239 13875 6245
rect 13817 6205 13829 6239
rect 13863 6236 13875 6239
rect 14336 6239 14372 6245
rect 14336 6236 14348 6239
rect 13863 6208 14348 6236
rect 13863 6205 13875 6208
rect 13817 6199 13875 6205
rect 14336 6205 14348 6208
rect 14336 6199 14372 6205
rect 14366 6196 14372 6199
rect 14424 6196 14430 6248
rect 9766 6128 9772 6180
rect 9824 6128 9830 6180
rect 14476 6168 14504 6412
rect 14918 6400 14924 6412
rect 14976 6400 14982 6452
rect 15010 6400 15016 6452
rect 15068 6440 15074 6452
rect 15473 6443 15531 6449
rect 15473 6440 15485 6443
rect 15068 6412 15485 6440
rect 15068 6400 15074 6412
rect 15473 6409 15485 6412
rect 15519 6440 15531 6443
rect 15562 6440 15568 6452
rect 15519 6412 15568 6440
rect 15519 6409 15531 6412
rect 15473 6403 15531 6409
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 16206 6440 16212 6452
rect 16167 6412 16212 6440
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 15102 6239 15160 6245
rect 15102 6205 15114 6239
rect 15148 6236 15160 6239
rect 15378 6236 15384 6248
rect 15148 6208 15384 6236
rect 15148 6205 15160 6208
rect 15102 6199 15160 6205
rect 15378 6196 15384 6208
rect 15436 6236 15442 6248
rect 15562 6236 15568 6248
rect 15436 6208 15568 6236
rect 15436 6196 15442 6208
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 16390 6236 16396 6248
rect 16351 6208 16396 6236
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 14292 6140 14504 6168
rect 10226 6100 10232 6112
rect 9048 6072 10232 6100
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10781 6103 10839 6109
rect 10781 6069 10793 6103
rect 10827 6100 10839 6103
rect 11514 6100 11520 6112
rect 10827 6072 11520 6100
rect 10827 6069 10839 6072
rect 10781 6063 10839 6069
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 12158 6060 12164 6112
rect 12216 6100 12222 6112
rect 12253 6103 12311 6109
rect 12253 6100 12265 6103
rect 12216 6072 12265 6100
rect 12216 6060 12222 6072
rect 12253 6069 12265 6072
rect 12299 6100 12311 6103
rect 14090 6100 14096 6112
rect 12299 6072 14096 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 14292 6109 14320 6140
rect 14277 6103 14335 6109
rect 14277 6069 14289 6103
rect 14323 6069 14335 6103
rect 14277 6063 14335 6069
rect 14366 6060 14372 6112
rect 14424 6100 14430 6112
rect 14461 6103 14519 6109
rect 14461 6100 14473 6103
rect 14424 6072 14473 6100
rect 14424 6060 14430 6072
rect 14461 6069 14473 6072
rect 14507 6069 14519 6103
rect 14461 6063 14519 6069
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 15105 6103 15163 6109
rect 15105 6100 15117 6103
rect 15068 6072 15117 6100
rect 15068 6060 15074 6072
rect 15105 6069 15117 6072
rect 15151 6069 15163 6103
rect 15105 6063 15163 6069
rect 1104 6010 17388 6032
rect 1104 5958 6410 6010
rect 6462 5958 6474 6010
rect 6526 5958 6538 6010
rect 6590 5958 6602 6010
rect 6654 5958 11838 6010
rect 11890 5958 11902 6010
rect 11954 5958 11966 6010
rect 12018 5958 12030 6010
rect 12082 5958 17388 6010
rect 1104 5936 17388 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 4249 5899 4307 5905
rect 4249 5896 4261 5899
rect 4212 5868 4261 5896
rect 4212 5856 4218 5868
rect 4249 5865 4261 5868
rect 4295 5865 4307 5899
rect 4249 5859 4307 5865
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5629 5899 5687 5905
rect 5629 5896 5641 5899
rect 4948 5868 5641 5896
rect 4948 5856 4954 5868
rect 5629 5865 5641 5868
rect 5675 5896 5687 5899
rect 5675 5868 7696 5896
rect 5675 5865 5687 5868
rect 5629 5859 5687 5865
rect 6914 5788 6920 5840
rect 6972 5788 6978 5840
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 4062 5720 4068 5772
rect 4120 5760 4126 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4120 5732 4445 5760
rect 4120 5720 4126 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 5810 5760 5816 5772
rect 5771 5732 5816 5760
rect 4433 5723 4491 5729
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 7374 5692 7380 5704
rect 7335 5664 7380 5692
rect 7374 5652 7380 5664
rect 7432 5652 7438 5704
rect 7668 5701 7696 5868
rect 10318 5856 10324 5908
rect 10376 5896 10382 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10376 5868 10701 5896
rect 10376 5856 10382 5868
rect 10689 5865 10701 5868
rect 10735 5865 10747 5899
rect 11514 5896 11520 5908
rect 10689 5859 10747 5865
rect 11440 5868 11520 5896
rect 8297 5831 8355 5837
rect 8297 5797 8309 5831
rect 8343 5828 8355 5831
rect 8662 5828 8668 5840
rect 8343 5800 8668 5828
rect 8343 5797 8355 5800
rect 8297 5791 8355 5797
rect 8662 5788 8668 5800
rect 8720 5788 8726 5840
rect 11440 5828 11468 5868
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 13817 5899 13875 5905
rect 13817 5865 13829 5899
rect 13863 5896 13875 5899
rect 15286 5896 15292 5908
rect 13863 5868 15292 5896
rect 13863 5865 13875 5868
rect 13817 5859 13875 5865
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 15620 5868 16681 5896
rect 15620 5856 15626 5868
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 16669 5859 16727 5865
rect 15194 5828 15200 5840
rect 11440 5800 12434 5828
rect 15155 5800 15200 5828
rect 10045 5763 10103 5769
rect 10045 5729 10057 5763
rect 10091 5760 10103 5763
rect 10594 5760 10600 5772
rect 10091 5732 10600 5760
rect 10091 5729 10103 5732
rect 10045 5723 10103 5729
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 10686 5720 10692 5772
rect 10744 5760 10750 5772
rect 10873 5763 10931 5769
rect 10873 5760 10885 5763
rect 10744 5732 10885 5760
rect 10744 5720 10750 5732
rect 10873 5729 10885 5732
rect 10919 5729 10931 5763
rect 10873 5723 10931 5729
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5692 7711 5695
rect 7742 5692 7748 5704
rect 7699 5664 7748 5692
rect 7699 5661 7711 5664
rect 7653 5655 7711 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 9861 5695 9919 5701
rect 9861 5692 9873 5695
rect 9824 5664 9873 5692
rect 9824 5652 9830 5664
rect 9861 5661 9873 5664
rect 9907 5661 9919 5695
rect 11440 5692 11468 5800
rect 11514 5763 11572 5769
rect 11514 5729 11526 5763
rect 11560 5760 11572 5763
rect 12406 5760 12434 5800
rect 15194 5788 15200 5800
rect 15252 5788 15258 5840
rect 16206 5788 16212 5840
rect 16264 5788 16270 5840
rect 12575 5763 12633 5769
rect 12575 5760 12587 5763
rect 11560 5732 12020 5760
rect 12406 5732 12587 5760
rect 11560 5729 11572 5732
rect 11514 5723 11572 5729
rect 11992 5701 12020 5732
rect 12575 5729 12587 5732
rect 12621 5729 12633 5763
rect 12710 5760 12716 5772
rect 12671 5732 12716 5760
rect 12575 5723 12633 5729
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 12802 5720 12808 5772
rect 12860 5760 12866 5772
rect 12989 5763 13047 5769
rect 12860 5732 12905 5760
rect 12860 5720 12866 5732
rect 12989 5729 13001 5763
rect 13035 5729 13047 5763
rect 12989 5723 13047 5729
rect 13633 5763 13691 5769
rect 13633 5729 13645 5763
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 11885 5695 11943 5701
rect 11885 5692 11897 5695
rect 11440 5664 11897 5692
rect 9861 5655 9919 5661
rect 11885 5661 11897 5664
rect 11931 5661 11943 5695
rect 11885 5655 11943 5661
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5692 12035 5695
rect 12728 5692 12756 5720
rect 12023 5664 12756 5692
rect 12023 5661 12035 5664
rect 11977 5655 12035 5661
rect 11054 5584 11060 5636
rect 11112 5624 11118 5636
rect 11333 5627 11391 5633
rect 11333 5624 11345 5627
rect 11112 5596 11345 5624
rect 11112 5584 11118 5596
rect 11333 5593 11345 5596
rect 11379 5624 11391 5627
rect 13004 5624 13032 5723
rect 11379 5596 13032 5624
rect 11379 5593 11391 5596
rect 11333 5587 11391 5593
rect 5902 5556 5908 5568
rect 5863 5528 5908 5556
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 8202 5556 8208 5568
rect 8163 5528 8208 5556
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 10229 5559 10287 5565
rect 10229 5525 10241 5559
rect 10275 5556 10287 5559
rect 10594 5556 10600 5568
rect 10275 5528 10600 5556
rect 10275 5525 10287 5528
rect 10229 5519 10287 5525
rect 10594 5516 10600 5528
rect 10652 5516 10658 5568
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 13648 5556 13676 5723
rect 14090 5652 14096 5704
rect 14148 5692 14154 5704
rect 14921 5695 14979 5701
rect 14921 5692 14933 5695
rect 14148 5664 14933 5692
rect 14148 5652 14154 5664
rect 14921 5661 14933 5664
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 15930 5556 15936 5568
rect 12492 5528 12537 5556
rect 13648 5528 15936 5556
rect 12492 5516 12498 5528
rect 15930 5516 15936 5528
rect 15988 5516 15994 5568
rect 1104 5466 17388 5488
rect 1104 5414 3696 5466
rect 3748 5414 3760 5466
rect 3812 5414 3824 5466
rect 3876 5414 3888 5466
rect 3940 5414 9124 5466
rect 9176 5414 9188 5466
rect 9240 5414 9252 5466
rect 9304 5414 9316 5466
rect 9368 5414 14552 5466
rect 14604 5414 14616 5466
rect 14668 5414 14680 5466
rect 14732 5414 14744 5466
rect 14796 5414 17388 5466
rect 1104 5392 17388 5414
rect 3510 5312 3516 5364
rect 3568 5352 3574 5364
rect 3697 5355 3755 5361
rect 3697 5352 3709 5355
rect 3568 5324 3709 5352
rect 3568 5312 3574 5324
rect 3697 5321 3709 5324
rect 3743 5321 3755 5355
rect 3697 5315 3755 5321
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 4522 5352 4528 5364
rect 4387 5324 4528 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 4522 5312 4528 5324
rect 4580 5352 4586 5364
rect 4798 5352 4804 5364
rect 4580 5324 4804 5352
rect 4580 5312 4586 5324
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5261 5355 5319 5361
rect 5261 5321 5273 5355
rect 5307 5352 5319 5355
rect 5442 5352 5448 5364
rect 5307 5324 5448 5352
rect 5307 5321 5319 5324
rect 5261 5315 5319 5321
rect 5442 5312 5448 5324
rect 5500 5352 5506 5364
rect 6086 5352 6092 5364
rect 5500 5324 6092 5352
rect 5500 5312 5506 5324
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 6825 5355 6883 5361
rect 6825 5321 6837 5355
rect 6871 5352 6883 5355
rect 7374 5352 7380 5364
rect 6871 5324 7380 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 11054 5352 11060 5364
rect 11015 5324 11060 5352
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 12768 5324 13829 5352
rect 12768 5312 12774 5324
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 13817 5315 13875 5321
rect 14366 5312 14372 5364
rect 14424 5312 14430 5364
rect 5718 5244 5724 5296
rect 5776 5284 5782 5296
rect 5776 5256 7236 5284
rect 5776 5244 5782 5256
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 5994 5216 6000 5228
rect 5859 5188 6000 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 5994 5176 6000 5188
rect 6052 5216 6058 5228
rect 6052 5188 7052 5216
rect 6052 5176 6058 5188
rect 1946 5148 1952 5160
rect 1907 5120 1952 5148
rect 1946 5108 1952 5120
rect 2004 5108 2010 5160
rect 4157 5151 4215 5157
rect 4157 5117 4169 5151
rect 4203 5148 4215 5151
rect 4338 5148 4344 5160
rect 4203 5120 4344 5148
rect 4203 5117 4215 5120
rect 4157 5111 4215 5117
rect 4338 5108 4344 5120
rect 4396 5108 4402 5160
rect 5442 5151 5500 5157
rect 5442 5117 5454 5151
rect 5488 5148 5500 5151
rect 5488 5120 5764 5148
rect 5488 5117 5500 5120
rect 5442 5111 5500 5117
rect 2222 5080 2228 5092
rect 2183 5052 2228 5080
rect 2222 5040 2228 5052
rect 2280 5040 2286 5092
rect 2958 5040 2964 5092
rect 3016 5040 3022 5092
rect 5736 5080 5764 5120
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 7024 5157 7052 5188
rect 7208 5157 7236 5256
rect 10226 5176 10232 5228
rect 10284 5216 10290 5228
rect 11238 5216 11244 5228
rect 10284 5188 11244 5216
rect 10284 5176 10290 5188
rect 11238 5176 11244 5188
rect 11296 5216 11302 5228
rect 12066 5216 12072 5228
rect 11296 5188 12072 5216
rect 11296 5176 11302 5188
rect 12066 5176 12072 5188
rect 12124 5176 12130 5228
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5216 12403 5219
rect 12434 5216 12440 5228
rect 12391 5188 12440 5216
rect 12391 5185 12403 5188
rect 12345 5179 12403 5185
rect 12434 5176 12440 5188
rect 12492 5176 12498 5228
rect 14090 5176 14096 5228
rect 14148 5216 14154 5228
rect 14277 5219 14335 5225
rect 14277 5216 14289 5219
rect 14148 5188 14289 5216
rect 14148 5176 14154 5188
rect 14277 5185 14289 5188
rect 14323 5185 14335 5219
rect 14384 5216 14412 5312
rect 14553 5219 14611 5225
rect 14553 5216 14565 5219
rect 14384 5188 14565 5216
rect 14277 5179 14335 5185
rect 14553 5185 14565 5188
rect 14599 5185 14611 5219
rect 14553 5179 14611 5185
rect 7009 5151 7067 5157
rect 5960 5120 6053 5148
rect 5960 5108 5966 5120
rect 7009 5117 7021 5151
rect 7055 5117 7067 5151
rect 7009 5111 7067 5117
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5117 7251 5151
rect 7193 5111 7251 5117
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 5920 5080 5948 5108
rect 7101 5083 7159 5089
rect 7101 5080 7113 5083
rect 5736 5052 7113 5080
rect 7101 5049 7113 5052
rect 7147 5049 7159 5083
rect 7101 5043 7159 5049
rect 5445 5015 5503 5021
rect 5445 4981 5457 5015
rect 5491 5012 5503 5015
rect 5994 5012 6000 5024
rect 5491 4984 6000 5012
rect 5491 4981 5503 4984
rect 5445 4975 5503 4981
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 7392 5012 7420 5111
rect 7742 5108 7748 5160
rect 7800 5148 7806 5160
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7800 5120 7941 5148
rect 7800 5108 7806 5120
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 10686 5151 10744 5157
rect 10686 5117 10698 5151
rect 10732 5117 10744 5151
rect 10686 5111 10744 5117
rect 11149 5151 11207 5157
rect 11149 5117 11161 5151
rect 11195 5117 11207 5151
rect 11149 5111 11207 5117
rect 8205 5083 8263 5089
rect 8205 5049 8217 5083
rect 8251 5080 8263 5083
rect 8478 5080 8484 5092
rect 8251 5052 8484 5080
rect 8251 5049 8263 5052
rect 8205 5043 8263 5049
rect 8478 5040 8484 5052
rect 8536 5040 8542 5092
rect 9490 5080 9496 5092
rect 9430 5052 9496 5080
rect 9490 5040 9496 5052
rect 9548 5040 9554 5092
rect 10701 5080 10729 5111
rect 11164 5080 11192 5111
rect 12618 5080 12624 5092
rect 10701 5052 12624 5080
rect 12618 5040 12624 5052
rect 12676 5040 12682 5092
rect 13354 5040 13360 5092
rect 13412 5040 13418 5092
rect 15010 5040 15016 5092
rect 15068 5040 15074 5092
rect 9674 5012 9680 5024
rect 6144 4984 7420 5012
rect 9635 4984 9680 5012
rect 6144 4972 6150 4984
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 10502 5012 10508 5024
rect 10463 4984 10508 5012
rect 10502 4972 10508 4984
rect 10560 4972 10566 5024
rect 10689 5015 10747 5021
rect 10689 4981 10701 5015
rect 10735 5012 10747 5015
rect 11054 5012 11060 5024
rect 10735 4984 11060 5012
rect 10735 4981 10747 4984
rect 10689 4975 10747 4981
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 16022 5012 16028 5024
rect 15983 4984 16028 5012
rect 16022 4972 16028 4984
rect 16080 4972 16086 5024
rect 1104 4922 17388 4944
rect 1104 4870 6410 4922
rect 6462 4870 6474 4922
rect 6526 4870 6538 4922
rect 6590 4870 6602 4922
rect 6654 4870 11838 4922
rect 11890 4870 11902 4922
rect 11954 4870 11966 4922
rect 12018 4870 12030 4922
rect 12082 4870 17388 4922
rect 1104 4848 17388 4870
rect 2958 4808 2964 4820
rect 2919 4780 2964 4808
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 4890 4808 4896 4820
rect 4264 4780 4896 4808
rect 2774 4632 2780 4684
rect 2832 4672 2838 4684
rect 4062 4672 4068 4684
rect 2832 4644 4068 4672
rect 2832 4632 2838 4644
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 4264 4681 4292 4780
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5994 4808 6000 4820
rect 5955 4780 6000 4808
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 9490 4808 9496 4820
rect 9451 4780 9496 4808
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 12802 4808 12808 4820
rect 12763 4780 12808 4808
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 13265 4811 13323 4817
rect 13265 4777 13277 4811
rect 13311 4808 13323 4811
rect 13354 4808 13360 4820
rect 13311 4780 13360 4808
rect 13311 4777 13323 4780
rect 13265 4771 13323 4777
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 14921 4811 14979 4817
rect 14921 4777 14933 4811
rect 14967 4808 14979 4811
rect 15010 4808 15016 4820
rect 14967 4780 15016 4808
rect 14967 4777 14979 4780
rect 14921 4771 14979 4777
rect 15010 4768 15016 4780
rect 15068 4768 15074 4820
rect 16206 4808 16212 4820
rect 16167 4780 16212 4808
rect 16206 4768 16212 4780
rect 16264 4768 16270 4820
rect 9766 4740 9772 4752
rect 7024 4712 9772 4740
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4641 4307 4675
rect 4249 4635 4307 4641
rect 1946 4564 1952 4616
rect 2004 4604 2010 4616
rect 4264 4604 4292 4635
rect 5626 4632 5632 4684
rect 5684 4632 5690 4684
rect 4522 4604 4528 4616
rect 2004 4576 4292 4604
rect 4483 4576 4528 4604
rect 2004 4564 2010 4576
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 7024 4604 7052 4712
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 10502 4740 10508 4752
rect 10463 4712 10508 4740
rect 10502 4700 10508 4712
rect 10560 4700 10566 4752
rect 12066 4740 12072 4752
rect 11730 4712 12072 4740
rect 12066 4700 12072 4712
rect 12124 4700 12130 4752
rect 15212 4712 16436 4740
rect 15212 4684 15240 4712
rect 16408 4684 16436 4712
rect 7098 4632 7104 4684
rect 7156 4672 7162 4684
rect 7193 4675 7251 4681
rect 7193 4672 7205 4675
rect 7156 4644 7205 4672
rect 7156 4632 7162 4644
rect 7193 4641 7205 4644
rect 7239 4672 7251 4675
rect 8386 4672 8392 4684
rect 7239 4644 8392 4672
rect 7239 4641 7251 4644
rect 7193 4635 7251 4641
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 8662 4672 8668 4684
rect 8619 4644 8668 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 10226 4672 10232 4684
rect 10187 4644 10232 4672
rect 9677 4635 9735 4641
rect 8294 4604 8300 4616
rect 4948 4576 7052 4604
rect 8255 4576 8300 4604
rect 4948 4564 4954 4576
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8018 4536 8024 4548
rect 5549 4508 8024 4536
rect 4062 4428 4068 4480
rect 4120 4468 4126 4480
rect 5549 4468 5577 4508
rect 8018 4496 8024 4508
rect 8076 4536 8082 4548
rect 9692 4536 9720 4635
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 12621 4675 12679 4681
rect 12621 4641 12633 4675
rect 12667 4641 12679 4675
rect 12621 4635 12679 4641
rect 9766 4564 9772 4616
rect 9824 4604 9830 4616
rect 12437 4607 12495 4613
rect 12437 4604 12449 4607
rect 9824 4576 12449 4604
rect 9824 4564 9830 4576
rect 12437 4573 12449 4576
rect 12483 4573 12495 4607
rect 12636 4604 12664 4635
rect 13354 4632 13360 4684
rect 13412 4672 13418 4684
rect 13449 4675 13507 4681
rect 13449 4672 13461 4675
rect 13412 4644 13461 4672
rect 13412 4632 13418 4644
rect 13449 4641 13461 4644
rect 13495 4641 13507 4675
rect 13449 4635 13507 4641
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 15194 4672 15200 4684
rect 14783 4644 15200 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 15194 4632 15200 4644
rect 15252 4632 15258 4684
rect 15746 4672 15752 4684
rect 15707 4644 15752 4672
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 16390 4672 16396 4684
rect 16303 4644 16396 4672
rect 16390 4632 16396 4644
rect 16448 4632 16454 4684
rect 13814 4604 13820 4616
rect 12636 4576 13820 4604
rect 12437 4567 12495 4573
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 8076 4508 9720 4536
rect 8076 4496 8082 4508
rect 4120 4440 5577 4468
rect 4120 4428 4126 4440
rect 6914 4428 6920 4480
rect 6972 4468 6978 4480
rect 7009 4471 7067 4477
rect 7009 4468 7021 4471
rect 6972 4440 7021 4468
rect 6972 4428 6978 4440
rect 7009 4437 7021 4440
rect 7055 4437 7067 4471
rect 7009 4431 7067 4437
rect 11977 4471 12035 4477
rect 11977 4437 11989 4471
rect 12023 4468 12035 4471
rect 12158 4468 12164 4480
rect 12023 4440 12164 4468
rect 12023 4437 12035 4440
rect 11977 4431 12035 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 15565 4471 15623 4477
rect 15565 4437 15577 4471
rect 15611 4468 15623 4471
rect 15654 4468 15660 4480
rect 15611 4440 15660 4468
rect 15611 4437 15623 4440
rect 15565 4431 15623 4437
rect 15654 4428 15660 4440
rect 15712 4428 15718 4480
rect 1104 4378 17388 4400
rect 1104 4326 3696 4378
rect 3748 4326 3760 4378
rect 3812 4326 3824 4378
rect 3876 4326 3888 4378
rect 3940 4326 9124 4378
rect 9176 4326 9188 4378
rect 9240 4326 9252 4378
rect 9304 4326 9316 4378
rect 9368 4326 14552 4378
rect 14604 4326 14616 4378
rect 14668 4326 14680 4378
rect 14732 4326 14744 4378
rect 14796 4326 17388 4378
rect 1104 4304 17388 4326
rect 5626 4264 5632 4276
rect 5587 4236 5632 4264
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 8018 4264 8024 4276
rect 7979 4236 8024 4264
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 10965 4267 11023 4273
rect 10965 4264 10977 4267
rect 8536 4236 10977 4264
rect 8536 4224 8542 4236
rect 10965 4233 10977 4236
rect 11011 4233 11023 4267
rect 12066 4264 12072 4276
rect 12027 4236 12072 4264
rect 10965 4227 11023 4233
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 15286 4224 15292 4276
rect 15344 4264 15350 4276
rect 15657 4267 15715 4273
rect 15657 4264 15669 4267
rect 15344 4236 15669 4264
rect 15344 4224 15350 4236
rect 15657 4233 15669 4236
rect 15703 4264 15715 4267
rect 16022 4264 16028 4276
rect 15703 4236 16028 4264
rect 15703 4233 15715 4236
rect 15657 4227 15715 4233
rect 16022 4224 16028 4236
rect 16080 4224 16086 4276
rect 4062 4156 4068 4208
rect 4120 4156 4126 4208
rect 6825 4199 6883 4205
rect 6825 4165 6837 4199
rect 6871 4165 6883 4199
rect 6825 4159 6883 4165
rect 4080 4128 4108 4156
rect 3252 4100 4108 4128
rect 3252 4069 3280 4100
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 6840 4128 6868 4159
rect 8386 4156 8392 4208
rect 8444 4196 8450 4208
rect 8665 4199 8723 4205
rect 8665 4196 8677 4199
rect 8444 4168 8677 4196
rect 8444 4156 8450 4168
rect 8665 4165 8677 4168
rect 8711 4165 8723 4199
rect 8665 4159 8723 4165
rect 8202 4128 8208 4140
rect 4212 4100 6868 4128
rect 6932 4100 8208 4128
rect 4212 4088 4218 4100
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4029 3295 4063
rect 3237 4023 3295 4029
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 3881 4063 3939 4069
rect 3881 4060 3893 4063
rect 3568 4032 3893 4060
rect 3568 4020 3574 4032
rect 3881 4029 3893 4032
rect 3927 4029 3939 4063
rect 3881 4023 3939 4029
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 4985 4063 5043 4069
rect 4985 4060 4997 4063
rect 4120 4032 4997 4060
rect 4120 4020 4126 4032
rect 4985 4029 4997 4032
rect 5031 4029 5043 4063
rect 5166 4060 5172 4072
rect 5127 4032 5172 4060
rect 4985 4023 5043 4029
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 6932 4060 6960 4100
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4128 9367 4131
rect 12526 4128 12532 4140
rect 9355 4100 10732 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 9692 4072 9720 4100
rect 5859 4032 6960 4060
rect 7009 4063 7067 4069
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 7009 4029 7021 4063
rect 7055 4029 7067 4063
rect 7009 4023 7067 4029
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4060 8171 4063
rect 8662 4060 8668 4072
rect 8159 4032 8668 4060
rect 8159 4029 8171 4032
rect 8113 4023 8171 4029
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 7024 3992 7052 4023
rect 8662 4020 8668 4032
rect 8720 4060 8726 4072
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 8720 4032 8861 4060
rect 8720 4020 8726 4032
rect 8849 4029 8861 4032
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 9401 4063 9459 4069
rect 9401 4029 9413 4063
rect 9447 4060 9459 4063
rect 9490 4060 9496 4072
rect 9447 4032 9496 4060
rect 9447 4029 9459 4032
rect 9401 4023 9459 4029
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 9772 4063 9830 4069
rect 9772 4060 9784 4063
rect 9732 4032 9784 4060
rect 9732 4020 9738 4032
rect 9772 4029 9784 4032
rect 9818 4029 9830 4063
rect 9772 4023 9830 4029
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 10008 4032 10425 4060
rect 10008 4020 10014 4032
rect 10413 4029 10425 4032
rect 10459 4029 10471 4063
rect 10594 4060 10600 4072
rect 10555 4032 10600 4060
rect 10413 4023 10471 4029
rect 10594 4020 10600 4032
rect 10652 4020 10658 4072
rect 10704 4069 10732 4100
rect 12406 4100 12532 4128
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4029 10747 4063
rect 10689 4023 10747 4029
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 12253 4063 12311 4069
rect 12253 4029 12265 4063
rect 12299 4060 12311 4063
rect 12406 4060 12434 4100
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 14090 4088 14096 4140
rect 14148 4128 14154 4140
rect 14461 4131 14519 4137
rect 14461 4128 14473 4131
rect 14148 4100 14473 4128
rect 14148 4088 14154 4100
rect 14461 4097 14473 4100
rect 14507 4128 14519 4131
rect 14918 4128 14924 4140
rect 14507 4100 14924 4128
rect 14507 4097 14519 4100
rect 14461 4091 14519 4097
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 12299 4032 12434 4060
rect 15286 4063 15344 4069
rect 12299 4029 12311 4032
rect 12253 4023 12311 4029
rect 15286 4029 15298 4063
rect 15332 4060 15344 4063
rect 15749 4063 15807 4069
rect 15749 4060 15761 4063
rect 15332 4032 15761 4060
rect 15332 4029 15344 4032
rect 15286 4023 15344 4029
rect 15749 4029 15761 4032
rect 15795 4060 15807 4063
rect 15838 4060 15844 4072
rect 15795 4032 15844 4060
rect 15795 4029 15807 4032
rect 15749 4023 15807 4029
rect 5592 3964 7052 3992
rect 9784 3964 10088 3992
rect 5592 3952 5598 3964
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 3421 3927 3479 3933
rect 3421 3924 3433 3927
rect 3384 3896 3433 3924
rect 3384 3884 3390 3896
rect 3421 3893 3433 3896
rect 3467 3893 3479 3927
rect 3421 3887 3479 3893
rect 4065 3927 4123 3933
rect 4065 3893 4077 3927
rect 4111 3924 4123 3927
rect 4706 3924 4712 3936
rect 4111 3896 4712 3924
rect 4111 3893 4123 3896
rect 4065 3887 4123 3893
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 4801 3927 4859 3933
rect 4801 3893 4813 3927
rect 4847 3924 4859 3927
rect 5718 3924 5724 3936
rect 4847 3896 5724 3924
rect 4847 3893 4859 3896
rect 4801 3887 4859 3893
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 5810 3884 5816 3936
rect 5868 3924 5874 3936
rect 8938 3924 8944 3936
rect 5868 3896 8944 3924
rect 5868 3884 5874 3896
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 9784 3933 9812 3964
rect 9769 3927 9827 3933
rect 9769 3924 9781 3927
rect 9548 3896 9781 3924
rect 9548 3884 9554 3896
rect 9769 3893 9781 3896
rect 9815 3893 9827 3927
rect 9950 3924 9956 3936
rect 9911 3896 9956 3924
rect 9769 3887 9827 3893
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10060 3924 10088 3964
rect 10796 3924 10824 4023
rect 15838 4020 15844 4032
rect 15896 4020 15902 4072
rect 16390 4069 16396 4072
rect 16385 4060 16396 4069
rect 16351 4032 16396 4060
rect 16385 4023 16396 4032
rect 16390 4020 16396 4023
rect 16448 4020 16454 4072
rect 13722 3952 13728 4004
rect 13780 3952 13786 4004
rect 14182 3992 14188 4004
rect 14143 3964 14188 3992
rect 14182 3952 14188 3964
rect 14240 3952 14246 4004
rect 12710 3924 12716 3936
rect 10060 3896 10824 3924
rect 12671 3896 12716 3924
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 15105 3927 15163 3933
rect 15105 3924 15117 3927
rect 15068 3896 15117 3924
rect 15068 3884 15074 3896
rect 15105 3893 15117 3896
rect 15151 3893 15163 3927
rect 15286 3924 15292 3936
rect 15247 3896 15292 3924
rect 15105 3887 15163 3893
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 16206 3924 16212 3936
rect 16167 3896 16212 3924
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 1104 3834 17388 3856
rect 1104 3782 6410 3834
rect 6462 3782 6474 3834
rect 6526 3782 6538 3834
rect 6590 3782 6602 3834
rect 6654 3782 11838 3834
rect 11890 3782 11902 3834
rect 11954 3782 11966 3834
rect 12018 3782 12030 3834
rect 12082 3782 17388 3834
rect 1104 3760 17388 3782
rect 2222 3680 2228 3732
rect 2280 3720 2286 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2280 3692 2697 3720
rect 2280 3680 2286 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3689 2927 3723
rect 2869 3683 2927 3689
rect 2884 3652 2912 3683
rect 4522 3680 4528 3732
rect 4580 3720 4586 3732
rect 4801 3723 4859 3729
rect 4801 3720 4813 3723
rect 4580 3692 4813 3720
rect 4580 3680 4586 3692
rect 4801 3689 4813 3692
rect 4847 3689 4859 3723
rect 4801 3683 4859 3689
rect 4985 3723 5043 3729
rect 4985 3689 4997 3723
rect 5031 3720 5043 3723
rect 5350 3720 5356 3732
rect 5031 3692 5356 3720
rect 5031 3689 5043 3692
rect 4985 3683 5043 3689
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 8570 3720 8576 3732
rect 5460 3692 8576 3720
rect 2792 3624 2912 3652
rect 2041 3587 2099 3593
rect 2041 3553 2053 3587
rect 2087 3553 2099 3587
rect 2041 3547 2099 3553
rect 2056 3448 2084 3547
rect 2792 3516 2820 3624
rect 3050 3612 3056 3664
rect 3108 3652 3114 3664
rect 5460 3652 5488 3692
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 9677 3723 9735 3729
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 9950 3720 9956 3732
rect 9723 3692 9956 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 10594 3720 10600 3732
rect 10152 3692 10600 3720
rect 3108 3624 5488 3652
rect 3108 3612 3114 3624
rect 6914 3612 6920 3664
rect 6972 3612 6978 3664
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 9582 3652 9588 3664
rect 8260 3624 9588 3652
rect 8260 3612 8266 3624
rect 9582 3612 9588 3624
rect 9640 3612 9646 3664
rect 10152 3652 10180 3692
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 10781 3723 10839 3729
rect 10781 3689 10793 3723
rect 10827 3720 10839 3723
rect 12986 3720 12992 3732
rect 10827 3692 12992 3720
rect 10827 3689 10839 3692
rect 10781 3683 10839 3689
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 13722 3720 13728 3732
rect 13683 3692 13728 3720
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 12526 3652 12532 3664
rect 9876 3624 10180 3652
rect 2866 3587 2924 3593
rect 2866 3553 2878 3587
rect 2912 3584 2924 3587
rect 4982 3587 5040 3593
rect 2912 3556 3372 3584
rect 2912 3553 2924 3556
rect 2866 3547 2924 3553
rect 3344 3525 3372 3556
rect 4982 3553 4994 3587
rect 5028 3584 5040 3587
rect 5028 3556 5488 3584
rect 5028 3553 5040 3556
rect 4982 3547 5040 3553
rect 3237 3519 3295 3525
rect 3237 3516 3249 3519
rect 2792 3488 3249 3516
rect 3237 3485 3249 3488
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 3329 3519 3387 3525
rect 3329 3485 3341 3519
rect 3375 3516 3387 3519
rect 3418 3516 3424 3528
rect 3375 3488 3424 3516
rect 3375 3485 3387 3488
rect 3329 3479 3387 3485
rect 3252 3448 3280 3479
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 5460 3525 5488 3556
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 8389 3587 8447 3593
rect 8389 3584 8401 3587
rect 8352 3556 8401 3584
rect 8352 3544 8358 3556
rect 8389 3553 8401 3556
rect 8435 3553 8447 3587
rect 8389 3547 8447 3553
rect 9674 3587 9732 3593
rect 9674 3553 9686 3587
rect 9720 3584 9732 3587
rect 9876 3584 9904 3624
rect 9720 3556 9904 3584
rect 9720 3553 9732 3556
rect 9674 3547 9732 3553
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3516 5503 3519
rect 5718 3516 5724 3528
rect 5491 3488 5724 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 7374 3516 7380 3528
rect 7335 3488 7380 3516
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 7653 3519 7711 3525
rect 7653 3485 7665 3519
rect 7699 3516 7711 3519
rect 7742 3516 7748 3528
rect 7699 3488 7748 3516
rect 7699 3485 7711 3488
rect 7653 3479 7711 3485
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 8404 3516 8432 3547
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 10152 3593 10180 3624
rect 10244 3624 12532 3652
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 10008 3556 10057 3584
rect 10008 3544 10014 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 8570 3516 8576 3528
rect 8404 3488 8576 3516
rect 8570 3476 8576 3488
rect 8628 3516 8634 3528
rect 10244 3516 10272 3624
rect 12526 3612 12532 3624
rect 12584 3652 12590 3664
rect 13354 3652 13360 3664
rect 12584 3624 13360 3652
rect 12584 3612 12590 3624
rect 13354 3612 13360 3624
rect 13412 3612 13418 3664
rect 15194 3652 15200 3664
rect 13556 3624 15200 3652
rect 10597 3587 10655 3593
rect 10597 3553 10609 3587
rect 10643 3553 10655 3587
rect 11422 3584 11428 3596
rect 11383 3556 11428 3584
rect 10597 3547 10655 3553
rect 8628 3488 10272 3516
rect 8628 3476 8634 3488
rect 4246 3448 4252 3460
rect 2056 3420 3188 3448
rect 3252 3420 4252 3448
rect 2225 3383 2283 3389
rect 2225 3349 2237 3383
rect 2271 3380 2283 3383
rect 3050 3380 3056 3392
rect 2271 3352 3056 3380
rect 2271 3349 2283 3352
rect 2225 3343 2283 3349
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 3160 3380 3188 3420
rect 4246 3408 4252 3420
rect 4304 3448 4310 3460
rect 4522 3448 4528 3460
rect 4304 3420 4528 3448
rect 4304 3408 4310 3420
rect 4522 3408 4528 3420
rect 4580 3408 4586 3460
rect 4632 3420 6132 3448
rect 4632 3380 4660 3420
rect 5350 3380 5356 3392
rect 3160 3352 4660 3380
rect 5311 3352 5356 3380
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 5905 3383 5963 3389
rect 5905 3349 5917 3383
rect 5951 3380 5963 3383
rect 5994 3380 6000 3392
rect 5951 3352 6000 3380
rect 5951 3349 5963 3352
rect 5905 3343 5963 3349
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 6104 3380 6132 3420
rect 8754 3408 8760 3460
rect 8812 3448 8818 3460
rect 10612 3448 10640 3547
rect 11422 3544 11428 3556
rect 11480 3544 11486 3596
rect 11606 3584 11612 3596
rect 11567 3556 11612 3584
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 11698 3544 11704 3596
rect 11756 3584 11762 3596
rect 11839 3587 11897 3593
rect 11756 3556 11801 3584
rect 11756 3544 11762 3556
rect 11839 3553 11851 3587
rect 11885 3584 11897 3587
rect 12158 3584 12164 3596
rect 11885 3556 12164 3584
rect 11885 3553 11897 3556
rect 11839 3547 11897 3553
rect 12158 3544 12164 3556
rect 12216 3544 12222 3596
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 13556 3593 13584 3624
rect 15194 3612 15200 3624
rect 15252 3612 15258 3664
rect 16206 3612 16212 3664
rect 16264 3612 16270 3664
rect 12621 3587 12679 3593
rect 12621 3584 12633 3587
rect 12492 3556 12633 3584
rect 12492 3544 12498 3556
rect 12621 3553 12633 3556
rect 12667 3553 12679 3587
rect 12621 3547 12679 3553
rect 13541 3587 13599 3593
rect 13541 3553 13553 3587
rect 13587 3553 13599 3587
rect 14918 3584 14924 3596
rect 14879 3556 14924 3584
rect 13541 3547 13599 3553
rect 13556 3516 13584 3547
rect 14918 3544 14924 3556
rect 14976 3544 14982 3596
rect 15194 3516 15200 3528
rect 8812 3420 10640 3448
rect 10701 3488 13584 3516
rect 15155 3488 15200 3516
rect 8812 3408 8818 3420
rect 7282 3380 7288 3392
rect 6104 3352 7288 3380
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 8202 3380 8208 3392
rect 8163 3352 8208 3380
rect 8202 3340 8208 3352
rect 8260 3340 8266 3392
rect 8478 3340 8484 3392
rect 8536 3380 8542 3392
rect 9493 3383 9551 3389
rect 9493 3380 9505 3383
rect 8536 3352 9505 3380
rect 8536 3340 8542 3352
rect 9493 3349 9505 3352
rect 9539 3349 9551 3383
rect 9493 3343 9551 3349
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 10701 3380 10729 3488
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 15838 3476 15844 3528
rect 15896 3516 15902 3528
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 15896 3488 16681 3516
rect 15896 3476 15902 3488
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 11977 3451 12035 3457
rect 11977 3417 11989 3451
rect 12023 3448 12035 3451
rect 13722 3448 13728 3460
rect 12023 3420 13728 3448
rect 12023 3417 12035 3420
rect 11977 3411 12035 3417
rect 13722 3408 13728 3420
rect 13780 3408 13786 3460
rect 9640 3352 10729 3380
rect 9640 3340 9646 3352
rect 11054 3340 11060 3392
rect 11112 3380 11118 3392
rect 12437 3383 12495 3389
rect 12437 3380 12449 3383
rect 11112 3352 12449 3380
rect 11112 3340 11118 3352
rect 12437 3349 12449 3352
rect 12483 3349 12495 3383
rect 12437 3343 12495 3349
rect 1104 3290 17388 3312
rect 1104 3238 3696 3290
rect 3748 3238 3760 3290
rect 3812 3238 3824 3290
rect 3876 3238 3888 3290
rect 3940 3238 9124 3290
rect 9176 3238 9188 3290
rect 9240 3238 9252 3290
rect 9304 3238 9316 3290
rect 9368 3238 14552 3290
rect 14604 3238 14616 3290
rect 14668 3238 14680 3290
rect 14732 3238 14744 3290
rect 14796 3238 17388 3290
rect 1104 3216 17388 3238
rect 1949 3179 2007 3185
rect 1949 3145 1961 3179
rect 1995 3176 2007 3179
rect 4062 3176 4068 3188
rect 1995 3148 4068 3176
rect 1995 3145 2007 3148
rect 1949 3139 2007 3145
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4522 3176 4528 3188
rect 4483 3148 4528 3176
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 7742 3136 7748 3188
rect 7800 3176 7806 3188
rect 9217 3179 9275 3185
rect 7800 3148 8800 3176
rect 7800 3136 7806 3148
rect 3970 3068 3976 3120
rect 4028 3108 4034 3120
rect 5810 3108 5816 3120
rect 4028 3080 5816 3108
rect 4028 3068 4034 3080
rect 5810 3068 5816 3080
rect 5868 3068 5874 3120
rect 1946 3000 1952 3052
rect 2004 3040 2010 3052
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 2004 3012 2329 3040
rect 2004 3000 2010 3012
rect 2317 3009 2329 3012
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 5123 3012 7021 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 474 2932 480 2984
rect 532 2972 538 2984
rect 1765 2975 1823 2981
rect 1765 2972 1777 2975
rect 532 2944 1777 2972
rect 532 2932 538 2944
rect 1765 2941 1777 2944
rect 1811 2941 1823 2975
rect 4080 2972 4108 3003
rect 4522 2972 4528 2984
rect 4080 2944 4528 2972
rect 1765 2935 1823 2941
rect 4522 2932 4528 2944
rect 4580 2972 4586 2984
rect 4650 2975 4708 2981
rect 4650 2972 4662 2975
rect 4580 2944 4662 2972
rect 4580 2932 4586 2944
rect 4650 2941 4662 2944
rect 4696 2972 4708 2975
rect 5169 2975 5227 2981
rect 5169 2972 5181 2975
rect 4696 2944 5181 2972
rect 4696 2941 4708 2944
rect 4650 2935 4708 2941
rect 5169 2941 5181 2944
rect 5215 2941 5227 2975
rect 5169 2935 5227 2941
rect 2593 2907 2651 2913
rect 2593 2873 2605 2907
rect 2639 2873 2651 2907
rect 2593 2867 2651 2873
rect 2608 2836 2636 2867
rect 3326 2864 3332 2916
rect 3384 2864 3390 2916
rect 5276 2904 5304 3012
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 8478 3040 8484 3052
rect 8439 3012 8484 3040
rect 7009 3003 7067 3009
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 8772 3049 8800 3148
rect 9217 3145 9229 3179
rect 9263 3176 9275 3179
rect 9490 3176 9496 3188
rect 9263 3148 9496 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 9490 3136 9496 3148
rect 9548 3136 9554 3188
rect 11422 3136 11428 3188
rect 11480 3176 11486 3188
rect 12069 3179 12127 3185
rect 12069 3176 12081 3179
rect 11480 3148 12081 3176
rect 11480 3136 11486 3148
rect 12069 3145 12081 3148
rect 12115 3145 12127 3179
rect 13814 3176 13820 3188
rect 13775 3148 13820 3176
rect 12069 3139 12127 3145
rect 13814 3136 13820 3148
rect 13872 3136 13878 3188
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 14461 3179 14519 3185
rect 14461 3176 14473 3179
rect 14240 3148 14473 3176
rect 14240 3136 14246 3148
rect 14461 3145 14473 3148
rect 14507 3145 14519 3179
rect 15010 3176 15016 3188
rect 14971 3148 15016 3176
rect 14461 3139 14519 3145
rect 15010 3136 15016 3148
rect 15068 3136 15074 3188
rect 15194 3136 15200 3188
rect 15252 3176 15258 3188
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 15252 3148 16129 3176
rect 15252 3136 15258 3148
rect 16117 3145 16129 3148
rect 16163 3145 16175 3179
rect 16117 3139 16175 3145
rect 15562 3108 15568 3120
rect 11348 3080 15568 3108
rect 8757 3043 8815 3049
rect 8757 3009 8769 3043
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3040 11023 3043
rect 11238 3040 11244 3052
rect 11011 3012 11244 3040
rect 11011 3009 11023 3012
rect 10965 3003 11023 3009
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 3896 2876 4660 2904
rect 3896 2836 3924 2876
rect 4632 2848 4660 2876
rect 4724 2876 5304 2904
rect 4724 2848 4752 2876
rect 5442 2864 5448 2916
rect 5500 2904 5506 2916
rect 5721 2907 5779 2913
rect 5721 2904 5733 2907
rect 5500 2876 5733 2904
rect 5500 2864 5506 2876
rect 5721 2873 5733 2876
rect 5767 2873 5779 2907
rect 8202 2904 8208 2916
rect 8050 2876 8208 2904
rect 5721 2867 5779 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 9674 2864 9680 2916
rect 9732 2864 9738 2916
rect 10594 2864 10600 2916
rect 10652 2904 10658 2916
rect 10689 2907 10747 2913
rect 10689 2904 10701 2907
rect 10652 2876 10701 2904
rect 10652 2864 10658 2876
rect 10689 2873 10701 2876
rect 10735 2873 10747 2907
rect 10689 2867 10747 2873
rect 2608 2808 3924 2836
rect 4614 2796 4620 2848
rect 4672 2796 4678 2848
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 4764 2808 4857 2836
rect 4764 2796 4770 2808
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 5813 2839 5871 2845
rect 5813 2836 5825 2839
rect 5224 2808 5825 2836
rect 5224 2796 5230 2808
rect 5813 2805 5825 2808
rect 5859 2836 5871 2839
rect 11348 2836 11376 3080
rect 15562 3068 15568 3080
rect 15620 3068 15626 3120
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 11756 3012 12725 3040
rect 11756 3000 11762 3012
rect 12268 2984 12296 3012
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 12713 3003 12771 3009
rect 15010 3000 15016 3052
rect 15068 3040 15074 3052
rect 15068 3012 15608 3040
rect 15068 3000 15074 3012
rect 12250 2972 12256 2984
rect 12163 2944 12256 2972
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 12621 2975 12679 2981
rect 12621 2972 12633 2975
rect 12406 2944 12633 2972
rect 5859 2808 11376 2836
rect 5859 2805 5871 2808
rect 5813 2799 5871 2805
rect 12158 2796 12164 2848
rect 12216 2836 12222 2848
rect 12253 2839 12311 2845
rect 12253 2836 12265 2839
rect 12216 2808 12265 2836
rect 12216 2796 12222 2808
rect 12253 2805 12265 2808
rect 12299 2836 12311 2839
rect 12406 2836 12434 2944
rect 12621 2941 12633 2944
rect 12667 2941 12679 2975
rect 13354 2972 13360 2984
rect 13315 2944 13360 2972
rect 12621 2935 12679 2941
rect 13354 2932 13360 2944
rect 13412 2932 13418 2984
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2972 14059 2975
rect 14274 2972 14280 2984
rect 14047 2944 14280 2972
rect 14047 2941 14059 2944
rect 14001 2935 14059 2941
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 15580 2981 15608 3012
rect 14642 2975 14700 2981
rect 14642 2941 14654 2975
rect 14688 2972 14700 2975
rect 15105 2975 15163 2981
rect 15105 2972 15117 2975
rect 14688 2944 15117 2972
rect 14688 2941 14700 2944
rect 14642 2935 14700 2941
rect 15105 2941 15117 2944
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 15565 2975 15623 2981
rect 15565 2941 15577 2975
rect 15611 2941 15623 2975
rect 15838 2972 15844 2984
rect 15799 2944 15844 2972
rect 15565 2935 15623 2941
rect 15120 2904 15148 2935
rect 15838 2932 15844 2944
rect 15896 2932 15902 2984
rect 15933 2975 15991 2981
rect 15933 2941 15945 2975
rect 15979 2972 15991 2975
rect 16022 2972 16028 2984
rect 15979 2944 16028 2972
rect 15979 2941 15991 2944
rect 15933 2935 15991 2941
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 15470 2904 15476 2916
rect 15120 2876 15476 2904
rect 15470 2864 15476 2876
rect 15528 2904 15534 2916
rect 15749 2907 15807 2913
rect 15749 2904 15761 2907
rect 15528 2876 15761 2904
rect 15528 2864 15534 2876
rect 15749 2873 15761 2876
rect 15795 2873 15807 2907
rect 15749 2867 15807 2873
rect 13170 2836 13176 2848
rect 12299 2808 12434 2836
rect 13131 2808 13176 2836
rect 12299 2805 12311 2808
rect 12253 2799 12311 2805
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 14645 2839 14703 2845
rect 14645 2805 14657 2839
rect 14691 2836 14703 2839
rect 15010 2836 15016 2848
rect 14691 2808 15016 2836
rect 14691 2805 14703 2808
rect 14645 2799 14703 2805
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 1104 2746 17388 2768
rect 1104 2694 6410 2746
rect 6462 2694 6474 2746
rect 6526 2694 6538 2746
rect 6590 2694 6602 2746
rect 6654 2694 11838 2746
rect 11890 2694 11902 2746
rect 11954 2694 11966 2746
rect 12018 2694 12030 2746
rect 12082 2694 17388 2746
rect 1104 2672 17388 2694
rect 2961 2635 3019 2641
rect 2961 2601 2973 2635
rect 3007 2632 3019 2635
rect 3418 2632 3424 2644
rect 3007 2604 3424 2632
rect 3007 2601 3019 2604
rect 2961 2595 3019 2601
rect 3418 2592 3424 2604
rect 3476 2632 3482 2644
rect 3476 2604 4292 2632
rect 3476 2592 3482 2604
rect 4154 2564 4160 2576
rect 3160 2536 4160 2564
rect 1854 2456 1860 2508
rect 1912 2496 1918 2508
rect 3160 2505 3188 2536
rect 4154 2524 4160 2536
rect 4212 2524 4218 2576
rect 4264 2564 4292 2604
rect 4614 2592 4620 2644
rect 4672 2632 4678 2644
rect 4801 2635 4859 2641
rect 4801 2632 4813 2635
rect 4672 2604 4813 2632
rect 4672 2592 4678 2604
rect 4801 2601 4813 2604
rect 4847 2601 4859 2635
rect 4801 2595 4859 2601
rect 5537 2635 5595 2641
rect 5537 2601 5549 2635
rect 5583 2632 5595 2635
rect 5626 2632 5632 2644
rect 5583 2604 5632 2632
rect 5583 2601 5595 2604
rect 5537 2595 5595 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 5994 2592 6000 2644
rect 6052 2632 6058 2644
rect 6052 2604 7236 2632
rect 6052 2592 6058 2604
rect 4522 2564 4528 2576
rect 4264 2536 4384 2564
rect 4483 2536 4528 2564
rect 1949 2499 2007 2505
rect 1949 2496 1961 2499
rect 1912 2468 1961 2496
rect 1912 2456 1918 2468
rect 1949 2465 1961 2468
rect 1995 2465 2007 2499
rect 1949 2459 2007 2465
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2465 3203 2499
rect 4246 2496 4252 2508
rect 4207 2468 4252 2496
rect 3145 2459 3203 2465
rect 4246 2456 4252 2468
rect 4304 2456 4310 2508
rect 4356 2496 4384 2536
rect 4522 2524 4528 2536
rect 4580 2524 4586 2576
rect 5718 2524 5724 2576
rect 5776 2564 5782 2576
rect 7208 2573 7236 2604
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 7432 2604 7481 2632
rect 7432 2592 7438 2604
rect 7469 2601 7481 2604
rect 7515 2601 7527 2635
rect 7469 2595 7527 2601
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 9674 2632 9680 2644
rect 8711 2604 9680 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 10505 2635 10563 2641
rect 10505 2601 10517 2635
rect 10551 2632 10563 2635
rect 10594 2632 10600 2644
rect 10551 2604 10600 2632
rect 10551 2601 10563 2604
rect 10505 2595 10563 2601
rect 10594 2592 10600 2604
rect 10652 2592 10658 2644
rect 10689 2635 10747 2641
rect 10689 2601 10701 2635
rect 10735 2632 10747 2635
rect 11422 2632 11428 2644
rect 10735 2604 11428 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 11422 2592 11428 2604
rect 11480 2592 11486 2644
rect 12250 2632 12256 2644
rect 12211 2604 12256 2632
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 15470 2632 15476 2644
rect 15431 2604 15476 2632
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 7101 2567 7159 2573
rect 7101 2564 7113 2567
rect 5776 2536 7113 2564
rect 5776 2524 5782 2536
rect 7101 2533 7113 2536
rect 7147 2533 7159 2567
rect 7101 2527 7159 2533
rect 7193 2567 7251 2573
rect 7193 2533 7205 2567
rect 7239 2533 7251 2567
rect 11054 2564 11060 2576
rect 7193 2527 7251 2533
rect 9876 2536 11060 2564
rect 4433 2499 4491 2505
rect 4433 2496 4445 2499
rect 4356 2468 4445 2496
rect 4433 2465 4445 2468
rect 4479 2465 4491 2499
rect 4433 2459 4491 2465
rect 4617 2499 4675 2505
rect 4617 2465 4629 2499
rect 4663 2496 4675 2499
rect 4706 2496 4712 2508
rect 4663 2468 4712 2496
rect 4663 2465 4675 2468
rect 4617 2459 4675 2465
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 5534 2499 5592 2505
rect 5534 2465 5546 2499
rect 5580 2496 5592 2499
rect 5994 2496 6000 2508
rect 5580 2468 6000 2496
rect 5580 2465 5592 2468
rect 5534 2459 5592 2465
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2496 8539 2499
rect 8570 2496 8576 2508
rect 8527 2468 8576 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2428 3387 2431
rect 4798 2428 4804 2440
rect 3375 2400 4804 2428
rect 3375 2397 3387 2400
rect 3329 2391 3387 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 5442 2428 5448 2440
rect 5184 2400 5448 2428
rect 2133 2363 2191 2369
rect 2133 2329 2145 2363
rect 2179 2360 2191 2363
rect 4338 2360 4344 2372
rect 2179 2332 4344 2360
rect 2179 2329 2191 2332
rect 2133 2323 2191 2329
rect 4338 2320 4344 2332
rect 4396 2360 4402 2372
rect 5184 2360 5212 2400
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 5350 2360 5356 2372
rect 4396 2332 5212 2360
rect 5263 2332 5356 2360
rect 4396 2320 4402 2332
rect 5350 2320 5356 2332
rect 5408 2360 5414 2372
rect 6932 2360 6960 2459
rect 5408 2332 6960 2360
rect 7300 2428 7328 2459
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 9876 2505 9904 2536
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 13170 2524 13176 2576
rect 13228 2524 13234 2576
rect 13722 2564 13728 2576
rect 13683 2536 13728 2564
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 15562 2524 15568 2576
rect 15620 2564 15626 2576
rect 15620 2536 15792 2564
rect 15620 2524 15626 2536
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2465 9919 2499
rect 9861 2459 9919 2465
rect 10045 2499 10103 2505
rect 10045 2465 10057 2499
rect 10091 2496 10103 2499
rect 10686 2499 10744 2505
rect 10686 2496 10698 2499
rect 10091 2468 10698 2496
rect 10091 2465 10103 2468
rect 10045 2459 10103 2465
rect 10686 2465 10698 2468
rect 10732 2496 10744 2499
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 10732 2468 11161 2496
rect 10732 2465 10744 2468
rect 10686 2459 10744 2465
rect 11149 2465 11161 2468
rect 11195 2496 11207 2499
rect 11606 2496 11612 2508
rect 11195 2468 11612 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 11606 2456 11612 2468
rect 11664 2456 11670 2508
rect 14001 2499 14059 2505
rect 14001 2465 14013 2499
rect 14047 2496 14059 2499
rect 14090 2496 14096 2508
rect 14047 2468 14096 2496
rect 14047 2465 14059 2468
rect 14001 2459 14059 2465
rect 14090 2456 14096 2468
rect 14148 2456 14154 2508
rect 15654 2496 15660 2508
rect 15615 2468 15660 2496
rect 15654 2456 15660 2468
rect 15712 2456 15718 2508
rect 15764 2505 15792 2536
rect 15749 2499 15807 2505
rect 15749 2465 15761 2499
rect 15795 2465 15807 2499
rect 15749 2459 15807 2465
rect 16669 2499 16727 2505
rect 16669 2465 16681 2499
rect 16715 2496 16727 2499
rect 17494 2496 17500 2508
rect 16715 2468 17500 2496
rect 16715 2465 16727 2468
rect 16669 2459 16727 2465
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 7300 2400 12434 2428
rect 5408 2320 5414 2332
rect 5626 2252 5632 2304
rect 5684 2292 5690 2304
rect 5905 2295 5963 2301
rect 5905 2292 5917 2295
rect 5684 2264 5917 2292
rect 5684 2252 5690 2264
rect 5905 2261 5917 2264
rect 5951 2292 5963 2295
rect 7300 2292 7328 2400
rect 11057 2363 11115 2369
rect 11057 2329 11069 2363
rect 11103 2360 11115 2363
rect 11422 2360 11428 2372
rect 11103 2332 11428 2360
rect 11103 2329 11115 2332
rect 11057 2323 11115 2329
rect 11422 2320 11428 2332
rect 11480 2320 11486 2372
rect 12406 2360 12434 2400
rect 12710 2360 12716 2372
rect 12406 2332 12716 2360
rect 12710 2320 12716 2332
rect 12768 2320 12774 2372
rect 16482 2292 16488 2304
rect 5951 2264 7328 2292
rect 16443 2264 16488 2292
rect 5951 2261 5963 2264
rect 5905 2255 5963 2261
rect 16482 2252 16488 2264
rect 16540 2252 16546 2304
rect 1104 2202 17388 2224
rect 1104 2150 3696 2202
rect 3748 2150 3760 2202
rect 3812 2150 3824 2202
rect 3876 2150 3888 2202
rect 3940 2150 9124 2202
rect 9176 2150 9188 2202
rect 9240 2150 9252 2202
rect 9304 2150 9316 2202
rect 9368 2150 14552 2202
rect 14604 2150 14616 2202
rect 14668 2150 14680 2202
rect 14732 2150 14744 2202
rect 14796 2150 17388 2202
rect 1104 2128 17388 2150
rect 4430 2048 4436 2100
rect 4488 2088 4494 2100
rect 16482 2088 16488 2100
rect 4488 2060 16488 2088
rect 4488 2048 4494 2060
rect 16482 2048 16488 2060
rect 16540 2048 16546 2100
<< via1 >>
rect 3696 18470 3748 18522
rect 3760 18470 3812 18522
rect 3824 18470 3876 18522
rect 3888 18470 3940 18522
rect 9124 18470 9176 18522
rect 9188 18470 9240 18522
rect 9252 18470 9304 18522
rect 9316 18470 9368 18522
rect 14552 18470 14604 18522
rect 14616 18470 14668 18522
rect 14680 18470 14732 18522
rect 14744 18470 14796 18522
rect 15292 18368 15344 18420
rect 7840 18343 7892 18352
rect 7840 18309 7849 18343
rect 7849 18309 7883 18343
rect 7883 18309 7892 18343
rect 7840 18300 7892 18309
rect 940 18232 992 18284
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 10140 18232 10192 18284
rect 4068 18164 4120 18216
rect 4804 18207 4856 18216
rect 4804 18173 4813 18207
rect 4813 18173 4847 18207
rect 4847 18173 4856 18207
rect 4804 18164 4856 18173
rect 5080 18164 5132 18216
rect 5540 18164 5592 18216
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 2320 18028 2372 18080
rect 4712 18028 4764 18080
rect 5264 18096 5316 18148
rect 8944 18164 8996 18216
rect 9864 18207 9916 18216
rect 9864 18173 9873 18207
rect 9873 18173 9907 18207
rect 9907 18173 9916 18207
rect 9864 18164 9916 18173
rect 16488 18300 16540 18352
rect 12164 18232 12216 18284
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 12900 18232 12952 18284
rect 15108 18207 15160 18216
rect 8576 18096 8628 18148
rect 11060 18096 11112 18148
rect 15108 18173 15117 18207
rect 15117 18173 15151 18207
rect 15151 18173 15160 18207
rect 15108 18164 15160 18173
rect 15292 18207 15344 18216
rect 15292 18173 15301 18207
rect 15301 18173 15335 18207
rect 15335 18173 15344 18207
rect 15292 18164 15344 18173
rect 15384 18164 15436 18216
rect 15200 18139 15252 18148
rect 15200 18105 15209 18139
rect 15209 18105 15243 18139
rect 15243 18105 15252 18139
rect 15200 18096 15252 18105
rect 6092 18028 6144 18080
rect 6828 18028 6880 18080
rect 12348 18028 12400 18080
rect 12900 18071 12952 18080
rect 12900 18037 12909 18071
rect 12909 18037 12943 18071
rect 12943 18037 12952 18071
rect 12900 18028 12952 18037
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 14924 18071 14976 18080
rect 14924 18037 14933 18071
rect 14933 18037 14967 18071
rect 14967 18037 14976 18071
rect 14924 18028 14976 18037
rect 15476 18028 15528 18080
rect 6410 17926 6462 17978
rect 6474 17926 6526 17978
rect 6538 17926 6590 17978
rect 6602 17926 6654 17978
rect 11838 17926 11890 17978
rect 11902 17926 11954 17978
rect 11966 17926 12018 17978
rect 12030 17926 12082 17978
rect 1952 17756 2004 17808
rect 6828 17824 6880 17876
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 15108 17867 15160 17876
rect 15108 17833 15117 17867
rect 15117 17833 15151 17867
rect 15151 17833 15160 17867
rect 15108 17824 15160 17833
rect 16488 17867 16540 17876
rect 16488 17833 16497 17867
rect 16497 17833 16531 17867
rect 16531 17833 16540 17867
rect 16488 17824 16540 17833
rect 6092 17799 6144 17808
rect 2320 17731 2372 17740
rect 2320 17697 2329 17731
rect 2329 17697 2363 17731
rect 2363 17697 2372 17731
rect 2320 17688 2372 17697
rect 6092 17765 6101 17799
rect 6101 17765 6135 17799
rect 6135 17765 6144 17799
rect 6092 17756 6144 17765
rect 8760 17756 8812 17808
rect 10048 17756 10100 17808
rect 13636 17756 13688 17808
rect 15200 17688 15252 17740
rect 17960 17688 18012 17740
rect 3516 17620 3568 17672
rect 5080 17620 5132 17672
rect 6736 17620 6788 17672
rect 7104 17663 7156 17672
rect 7104 17629 7113 17663
rect 7113 17629 7147 17663
rect 7147 17629 7156 17663
rect 7104 17620 7156 17629
rect 9772 17663 9824 17672
rect 2504 17527 2556 17536
rect 2504 17493 2513 17527
rect 2513 17493 2547 17527
rect 2547 17493 2556 17527
rect 2504 17484 2556 17493
rect 3332 17527 3384 17536
rect 3332 17493 3341 17527
rect 3341 17493 3375 17527
rect 3375 17493 3384 17527
rect 3332 17484 3384 17493
rect 4804 17484 4856 17536
rect 5356 17484 5408 17536
rect 9772 17629 9781 17663
rect 9781 17629 9815 17663
rect 9815 17629 9824 17663
rect 9772 17620 9824 17629
rect 12900 17620 12952 17672
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 15108 17552 15160 17604
rect 10876 17484 10928 17536
rect 12440 17484 12492 17536
rect 15384 17484 15436 17536
rect 3696 17382 3748 17434
rect 3760 17382 3812 17434
rect 3824 17382 3876 17434
rect 3888 17382 3940 17434
rect 9124 17382 9176 17434
rect 9188 17382 9240 17434
rect 9252 17382 9304 17434
rect 9316 17382 9368 17434
rect 14552 17382 14604 17434
rect 14616 17382 14668 17434
rect 14680 17382 14732 17434
rect 14744 17382 14796 17434
rect 3332 17280 3384 17332
rect 5080 17144 5132 17196
rect 2412 17076 2464 17128
rect 4804 17119 4856 17128
rect 4804 17085 4813 17119
rect 4813 17085 4847 17119
rect 4847 17085 4856 17119
rect 5264 17119 5316 17128
rect 4804 17076 4856 17085
rect 5264 17085 5273 17119
rect 5273 17085 5307 17119
rect 5307 17085 5316 17119
rect 5264 17076 5316 17085
rect 5356 17076 5408 17128
rect 7104 17280 7156 17332
rect 15568 17280 15620 17332
rect 6736 17212 6788 17264
rect 7656 17144 7708 17196
rect 10140 17144 10192 17196
rect 14924 17187 14976 17196
rect 14924 17153 14933 17187
rect 14933 17153 14967 17187
rect 14967 17153 14976 17187
rect 14924 17144 14976 17153
rect 7840 17076 7892 17128
rect 4436 17008 4488 17060
rect 4528 17051 4580 17060
rect 4528 17017 4537 17051
rect 4537 17017 4571 17051
rect 4571 17017 4580 17051
rect 5540 17051 5592 17060
rect 4528 17008 4580 17017
rect 5540 17017 5549 17051
rect 5549 17017 5583 17051
rect 5583 17017 5592 17051
rect 5540 17008 5592 17017
rect 8208 17051 8260 17060
rect 8208 17017 8217 17051
rect 8217 17017 8251 17051
rect 8251 17017 8260 17051
rect 8208 17008 8260 17017
rect 9496 17008 9548 17060
rect 2872 16940 2924 16992
rect 3240 16940 3292 16992
rect 5172 16940 5224 16992
rect 7656 16940 7708 16992
rect 7932 16940 7984 16992
rect 10508 16983 10560 16992
rect 10508 16949 10517 16983
rect 10517 16949 10551 16983
rect 10551 16949 10560 16983
rect 10508 16940 10560 16949
rect 12256 16983 12308 16992
rect 12256 16949 12265 16983
rect 12265 16949 12299 16983
rect 12299 16949 12308 16983
rect 12256 16940 12308 16949
rect 14096 17076 14148 17128
rect 13176 17008 13228 17060
rect 13728 17051 13780 17060
rect 13728 17017 13737 17051
rect 13737 17017 13771 17051
rect 13771 17017 13780 17051
rect 13728 17008 13780 17017
rect 15936 17008 15988 17060
rect 15292 16940 15344 16992
rect 6410 16838 6462 16890
rect 6474 16838 6526 16890
rect 6538 16838 6590 16890
rect 6602 16838 6654 16890
rect 11838 16838 11890 16890
rect 11902 16838 11954 16890
rect 11966 16838 12018 16890
rect 12030 16838 12082 16890
rect 3332 16736 3384 16788
rect 7196 16736 7248 16788
rect 8208 16779 8260 16788
rect 8208 16745 8217 16779
rect 8217 16745 8251 16779
rect 8251 16745 8260 16779
rect 8208 16736 8260 16745
rect 9772 16736 9824 16788
rect 10416 16736 10468 16788
rect 12440 16736 12492 16788
rect 13176 16779 13228 16788
rect 13176 16745 13185 16779
rect 13185 16745 13219 16779
rect 13219 16745 13228 16779
rect 13176 16736 13228 16745
rect 13636 16779 13688 16788
rect 13636 16745 13645 16779
rect 13645 16745 13679 16779
rect 13679 16745 13688 16779
rect 13636 16736 13688 16745
rect 5172 16711 5224 16720
rect 5172 16677 5181 16711
rect 5181 16677 5215 16711
rect 5215 16677 5224 16711
rect 5172 16668 5224 16677
rect 5908 16668 5960 16720
rect 7932 16711 7984 16720
rect 7932 16677 7941 16711
rect 7941 16677 7975 16711
rect 7975 16677 7984 16711
rect 7932 16668 7984 16677
rect 4160 16600 4212 16652
rect 4804 16600 4856 16652
rect 7656 16643 7708 16652
rect 7656 16609 7665 16643
rect 7665 16609 7699 16643
rect 7699 16609 7708 16643
rect 7656 16600 7708 16609
rect 7840 16643 7892 16652
rect 7840 16609 7849 16643
rect 7849 16609 7883 16643
rect 7883 16609 7892 16643
rect 7840 16600 7892 16609
rect 8208 16600 8260 16652
rect 9956 16600 10008 16652
rect 10508 16600 10560 16652
rect 10692 16600 10744 16652
rect 13360 16668 13412 16720
rect 12256 16600 12308 16652
rect 13268 16600 13320 16652
rect 15384 16736 15436 16788
rect 15936 16779 15988 16788
rect 15936 16745 15945 16779
rect 15945 16745 15979 16779
rect 15979 16745 15988 16779
rect 15936 16736 15988 16745
rect 3240 16575 3292 16584
rect 3240 16541 3249 16575
rect 3249 16541 3283 16575
rect 3283 16541 3292 16575
rect 3240 16532 3292 16541
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 12440 16532 12492 16541
rect 1492 16464 1544 16516
rect 2596 16439 2648 16448
rect 2596 16405 2605 16439
rect 2605 16405 2639 16439
rect 2639 16405 2648 16439
rect 2596 16396 2648 16405
rect 3332 16396 3384 16448
rect 12072 16464 12124 16516
rect 12348 16464 12400 16516
rect 15200 16643 15252 16652
rect 15200 16609 15212 16643
rect 15212 16609 15246 16643
rect 15246 16609 15252 16643
rect 16120 16643 16172 16652
rect 15200 16600 15252 16609
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 16120 16464 16172 16516
rect 10140 16396 10192 16448
rect 10416 16396 10468 16448
rect 15200 16396 15252 16448
rect 3696 16294 3748 16346
rect 3760 16294 3812 16346
rect 3824 16294 3876 16346
rect 3888 16294 3940 16346
rect 9124 16294 9176 16346
rect 9188 16294 9240 16346
rect 9252 16294 9304 16346
rect 9316 16294 9368 16346
rect 14552 16294 14604 16346
rect 14616 16294 14668 16346
rect 14680 16294 14732 16346
rect 14744 16294 14796 16346
rect 2596 16192 2648 16244
rect 4436 16235 4488 16244
rect 1492 16099 1544 16108
rect 1492 16065 1501 16099
rect 1501 16065 1535 16099
rect 1535 16065 1544 16099
rect 1492 16056 1544 16065
rect 2504 16056 2556 16108
rect 1676 16031 1728 16040
rect 1676 15997 1685 16031
rect 1685 15997 1719 16031
rect 1719 15997 1728 16031
rect 1676 15988 1728 15997
rect 3332 15988 3384 16040
rect 3240 15920 3292 15972
rect 4436 16201 4445 16235
rect 4445 16201 4479 16235
rect 4479 16201 4488 16235
rect 4436 16192 4488 16201
rect 5908 16235 5960 16244
rect 5908 16201 5917 16235
rect 5917 16201 5951 16235
rect 5951 16201 5960 16235
rect 5908 16192 5960 16201
rect 7656 16235 7708 16244
rect 7656 16201 7665 16235
rect 7665 16201 7699 16235
rect 7699 16201 7708 16235
rect 7656 16192 7708 16201
rect 8760 16235 8812 16244
rect 8760 16201 8769 16235
rect 8769 16201 8803 16235
rect 8803 16201 8812 16235
rect 8760 16192 8812 16201
rect 9496 16192 9548 16244
rect 13728 16192 13780 16244
rect 15292 16235 15344 16244
rect 15292 16201 15301 16235
rect 15301 16201 15335 16235
rect 15335 16201 15344 16235
rect 15292 16192 15344 16201
rect 9864 16124 9916 16176
rect 7932 16056 7984 16108
rect 4620 16031 4672 16040
rect 4620 15997 4629 16031
rect 4629 15997 4663 16031
rect 4663 15997 4672 16031
rect 4620 15988 4672 15997
rect 8208 16031 8260 16040
rect 4436 15920 4488 15972
rect 2044 15852 2096 15904
rect 2596 15852 2648 15904
rect 4528 15852 4580 15904
rect 8208 15997 8217 16031
rect 8217 15997 8251 16031
rect 8251 15997 8260 16031
rect 8208 15988 8260 15997
rect 8944 16031 8996 16040
rect 8944 15997 8953 16031
rect 8953 15997 8987 16031
rect 8987 15997 8996 16031
rect 8944 15988 8996 15997
rect 9680 15920 9732 15972
rect 7104 15852 7156 15904
rect 8208 15852 8260 15904
rect 9864 15852 9916 15904
rect 10416 15895 10468 15904
rect 10416 15861 10425 15895
rect 10425 15861 10459 15895
rect 10459 15861 10468 15895
rect 10416 15852 10468 15861
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 11244 15988 11296 16040
rect 12072 16031 12124 16040
rect 12072 15997 12081 16031
rect 12081 15997 12115 16031
rect 12115 15997 12124 16031
rect 12072 15988 12124 15997
rect 12164 15988 12216 16040
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 13268 16031 13320 16040
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 13912 16031 13964 16040
rect 13912 15997 13921 16031
rect 13921 15997 13955 16031
rect 13955 15997 13964 16031
rect 13912 15988 13964 15997
rect 15016 15988 15068 16040
rect 16580 16056 16632 16108
rect 16120 15988 16172 16040
rect 12348 15963 12400 15972
rect 12348 15929 12357 15963
rect 12357 15929 12391 15963
rect 12391 15929 12400 15963
rect 12348 15920 12400 15929
rect 14096 15963 14148 15972
rect 14096 15929 14105 15963
rect 14105 15929 14139 15963
rect 14139 15929 14148 15963
rect 14096 15920 14148 15929
rect 14924 15920 14976 15972
rect 10600 15852 10652 15861
rect 12716 15852 12768 15904
rect 14280 15852 14332 15904
rect 16212 15852 16264 15904
rect 6410 15750 6462 15802
rect 6474 15750 6526 15802
rect 6538 15750 6590 15802
rect 6602 15750 6654 15802
rect 11838 15750 11890 15802
rect 11902 15750 11954 15802
rect 11966 15750 12018 15802
rect 12030 15750 12082 15802
rect 5540 15648 5592 15700
rect 9956 15580 10008 15632
rect 11244 15648 11296 15700
rect 13268 15691 13320 15700
rect 13268 15657 13277 15691
rect 13277 15657 13311 15691
rect 13311 15657 13320 15691
rect 13268 15648 13320 15657
rect 12716 15580 12768 15632
rect 15200 15623 15252 15632
rect 15200 15589 15209 15623
rect 15209 15589 15243 15623
rect 15243 15589 15252 15623
rect 15200 15580 15252 15589
rect 16212 15580 16264 15632
rect 2964 15512 3016 15564
rect 4620 15512 4672 15564
rect 6000 15512 6052 15564
rect 6828 15512 6880 15564
rect 7104 15512 7156 15564
rect 8116 15555 8168 15564
rect 2228 15444 2280 15496
rect 8116 15521 8125 15555
rect 8125 15521 8159 15555
rect 8159 15521 8168 15555
rect 8116 15512 8168 15521
rect 9864 15555 9916 15564
rect 9864 15521 9873 15555
rect 9873 15521 9907 15555
rect 9907 15521 9916 15555
rect 9864 15512 9916 15521
rect 10600 15512 10652 15564
rect 10876 15555 10928 15564
rect 10876 15521 10885 15555
rect 10885 15521 10919 15555
rect 10919 15521 10928 15555
rect 10876 15512 10928 15521
rect 13360 15512 13412 15564
rect 11244 15444 11296 15496
rect 14004 15444 14056 15496
rect 1860 15351 1912 15360
rect 1860 15317 1869 15351
rect 1869 15317 1903 15351
rect 1903 15317 1912 15351
rect 1860 15308 1912 15317
rect 4620 15351 4672 15360
rect 4620 15317 4629 15351
rect 4629 15317 4663 15351
rect 4663 15317 4672 15351
rect 4620 15308 4672 15317
rect 6736 15308 6788 15360
rect 7564 15308 7616 15360
rect 15016 15308 15068 15360
rect 3696 15206 3748 15258
rect 3760 15206 3812 15258
rect 3824 15206 3876 15258
rect 3888 15206 3940 15258
rect 9124 15206 9176 15258
rect 9188 15206 9240 15258
rect 9252 15206 9304 15258
rect 9316 15206 9368 15258
rect 14552 15206 14604 15258
rect 14616 15206 14668 15258
rect 14680 15206 14732 15258
rect 14744 15206 14796 15258
rect 1676 15104 1728 15156
rect 4160 15104 4212 15156
rect 6736 15104 6788 15156
rect 5540 15036 5592 15088
rect 8208 15104 8260 15156
rect 10600 15104 10652 15156
rect 10876 15104 10928 15156
rect 1952 14943 2004 14952
rect 1952 14909 1961 14943
rect 1961 14909 1995 14943
rect 1995 14909 2004 14943
rect 1952 14900 2004 14909
rect 3976 14943 4028 14952
rect 3976 14909 3985 14943
rect 3985 14909 4019 14943
rect 4019 14909 4028 14943
rect 3976 14900 4028 14909
rect 4344 14900 4396 14952
rect 5816 14943 5868 14952
rect 5816 14909 5825 14943
rect 5825 14909 5859 14943
rect 5859 14909 5868 14943
rect 5816 14900 5868 14909
rect 9680 14968 9732 15020
rect 10876 14968 10928 15020
rect 6736 14900 6788 14952
rect 11336 14943 11388 14952
rect 11336 14909 11345 14943
rect 11345 14909 11379 14943
rect 11379 14909 11388 14943
rect 11336 14900 11388 14909
rect 3700 14875 3752 14884
rect 2228 14807 2280 14816
rect 2228 14773 2237 14807
rect 2237 14773 2271 14807
rect 2271 14773 2280 14807
rect 2228 14764 2280 14773
rect 3700 14841 3709 14875
rect 3709 14841 3743 14875
rect 3743 14841 3752 14875
rect 3700 14832 3752 14841
rect 5724 14832 5776 14884
rect 7564 14832 7616 14884
rect 5816 14764 5868 14816
rect 6000 14764 6052 14816
rect 9772 14832 9824 14884
rect 14096 15104 14148 15156
rect 13820 15036 13872 15088
rect 12808 14900 12860 14952
rect 14188 14968 14240 15020
rect 14832 14968 14884 15020
rect 15476 14968 15528 15020
rect 13820 14943 13872 14952
rect 12992 14832 13044 14884
rect 13820 14909 13829 14943
rect 13829 14909 13863 14943
rect 13863 14909 13872 14943
rect 13820 14900 13872 14909
rect 16396 14943 16448 14952
rect 16396 14909 16405 14943
rect 16405 14909 16439 14943
rect 16439 14909 16448 14943
rect 16396 14900 16448 14909
rect 13176 14764 13228 14816
rect 13820 14764 13872 14816
rect 14004 14764 14056 14816
rect 14372 14832 14424 14884
rect 14832 14764 14884 14816
rect 14924 14764 14976 14816
rect 16120 14764 16172 14816
rect 6410 14662 6462 14714
rect 6474 14662 6526 14714
rect 6538 14662 6590 14714
rect 6602 14662 6654 14714
rect 11838 14662 11890 14714
rect 11902 14662 11954 14714
rect 11966 14662 12018 14714
rect 12030 14662 12082 14714
rect 1860 14560 1912 14612
rect 3700 14560 3752 14612
rect 5816 14560 5868 14612
rect 2044 14424 2096 14476
rect 2228 14492 2280 14544
rect 4436 14492 4488 14544
rect 4620 14492 4672 14544
rect 6736 14535 6788 14544
rect 6736 14501 6745 14535
rect 6745 14501 6779 14535
rect 6779 14501 6788 14535
rect 6736 14492 6788 14501
rect 2964 14467 3016 14476
rect 2964 14433 2973 14467
rect 2973 14433 3007 14467
rect 3007 14433 3016 14467
rect 2964 14424 3016 14433
rect 3976 14424 4028 14476
rect 6644 14467 6696 14476
rect 5540 14356 5592 14408
rect 6644 14433 6653 14467
rect 6653 14433 6687 14467
rect 6687 14433 6696 14467
rect 6644 14424 6696 14433
rect 8944 14560 8996 14612
rect 9772 14560 9824 14612
rect 13912 14560 13964 14612
rect 15016 14560 15068 14612
rect 8116 14492 8168 14544
rect 10692 14492 10744 14544
rect 12164 14492 12216 14544
rect 13176 14492 13228 14544
rect 9496 14467 9548 14476
rect 9496 14433 9505 14467
rect 9505 14433 9539 14467
rect 9539 14433 9548 14467
rect 9496 14424 9548 14433
rect 10876 14424 10928 14476
rect 14464 14424 14516 14476
rect 14924 14467 14976 14476
rect 14924 14433 14930 14467
rect 14930 14433 14964 14467
rect 14964 14433 14976 14467
rect 14924 14424 14976 14433
rect 13084 14356 13136 14408
rect 15016 14356 15068 14408
rect 8944 14288 8996 14340
rect 10600 14288 10652 14340
rect 12808 14288 12860 14340
rect 6000 14220 6052 14272
rect 7012 14263 7064 14272
rect 7012 14229 7021 14263
rect 7021 14229 7055 14263
rect 7055 14229 7064 14263
rect 7012 14220 7064 14229
rect 12900 14263 12952 14272
rect 12900 14229 12909 14263
rect 12909 14229 12943 14263
rect 12943 14229 12952 14263
rect 12900 14220 12952 14229
rect 13636 14263 13688 14272
rect 13636 14229 13645 14263
rect 13645 14229 13679 14263
rect 13679 14229 13688 14263
rect 13636 14220 13688 14229
rect 16212 14220 16264 14272
rect 3696 14118 3748 14170
rect 3760 14118 3812 14170
rect 3824 14118 3876 14170
rect 3888 14118 3940 14170
rect 9124 14118 9176 14170
rect 9188 14118 9240 14170
rect 9252 14118 9304 14170
rect 9316 14118 9368 14170
rect 14552 14118 14604 14170
rect 14616 14118 14668 14170
rect 14680 14118 14732 14170
rect 14744 14118 14796 14170
rect 5540 14016 5592 14068
rect 5724 14059 5776 14068
rect 5724 14025 5733 14059
rect 5733 14025 5767 14059
rect 5767 14025 5776 14059
rect 5724 14016 5776 14025
rect 6736 14016 6788 14068
rect 3516 13991 3568 14000
rect 3516 13957 3525 13991
rect 3525 13957 3559 13991
rect 3559 13957 3568 13991
rect 3516 13948 3568 13957
rect 4160 13880 4212 13932
rect 4344 13948 4396 14000
rect 9496 14016 9548 14068
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 12164 14016 12216 14068
rect 13084 14059 13136 14068
rect 13084 14025 13093 14059
rect 13093 14025 13127 14059
rect 13127 14025 13136 14059
rect 13084 14016 13136 14025
rect 13268 14016 13320 14068
rect 13912 14016 13964 14068
rect 14372 14016 14424 14068
rect 7012 13880 7064 13932
rect 9680 13948 9732 14000
rect 9588 13880 9640 13932
rect 3516 13812 3568 13864
rect 4436 13855 4488 13864
rect 4436 13821 4445 13855
rect 4445 13821 4479 13855
rect 4479 13821 4488 13855
rect 4436 13812 4488 13821
rect 6644 13812 6696 13864
rect 8760 13812 8812 13864
rect 8944 13812 8996 13864
rect 11152 13855 11204 13864
rect 11152 13821 11161 13855
rect 11161 13821 11195 13855
rect 11195 13821 11204 13855
rect 11152 13812 11204 13821
rect 13820 13948 13872 14000
rect 15384 13948 15436 14000
rect 14096 13880 14148 13932
rect 13820 13812 13872 13864
rect 15108 13812 15160 13864
rect 16304 13855 16356 13864
rect 16304 13821 16313 13855
rect 16313 13821 16347 13855
rect 16347 13821 16356 13855
rect 16304 13812 16356 13821
rect 7288 13744 7340 13796
rect 10600 13744 10652 13796
rect 13360 13744 13412 13796
rect 2688 13719 2740 13728
rect 2688 13685 2697 13719
rect 2697 13685 2731 13719
rect 2731 13685 2740 13719
rect 2688 13676 2740 13685
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 10416 13676 10468 13728
rect 11336 13719 11388 13728
rect 11336 13685 11345 13719
rect 11345 13685 11379 13719
rect 11379 13685 11388 13719
rect 11336 13676 11388 13685
rect 13268 13719 13320 13728
rect 13268 13685 13277 13719
rect 13277 13685 13311 13719
rect 13311 13685 13320 13719
rect 13268 13676 13320 13685
rect 16028 13676 16080 13728
rect 6410 13574 6462 13626
rect 6474 13574 6526 13626
rect 6538 13574 6590 13626
rect 6602 13574 6654 13626
rect 11838 13574 11890 13626
rect 11902 13574 11954 13626
rect 11966 13574 12018 13626
rect 12030 13574 12082 13626
rect 2964 13472 3016 13524
rect 7288 13472 7340 13524
rect 10048 13472 10100 13524
rect 1400 13404 1452 13456
rect 2688 13404 2740 13456
rect 5540 13404 5592 13456
rect 13636 13472 13688 13524
rect 16488 13472 16540 13524
rect 4988 13379 5040 13388
rect 4988 13345 4997 13379
rect 4997 13345 5031 13379
rect 5031 13345 5040 13379
rect 4988 13336 5040 13345
rect 5172 13379 5224 13388
rect 5172 13345 5181 13379
rect 5181 13345 5215 13379
rect 5215 13345 5224 13379
rect 5172 13336 5224 13345
rect 5264 13268 5316 13320
rect 7104 13336 7156 13388
rect 11704 13404 11756 13456
rect 10600 13379 10652 13388
rect 7564 13268 7616 13320
rect 10600 13345 10609 13379
rect 10609 13345 10643 13379
rect 10643 13345 10652 13379
rect 10600 13336 10652 13345
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 12992 13336 13044 13345
rect 13360 13336 13412 13388
rect 16396 13336 16448 13388
rect 7932 13268 7984 13320
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 7840 13200 7892 13252
rect 11152 13200 11204 13252
rect 13820 13243 13872 13252
rect 13820 13209 13829 13243
rect 13829 13209 13863 13243
rect 13863 13209 13872 13243
rect 13820 13200 13872 13209
rect 15200 13200 15252 13252
rect 16304 13200 16356 13252
rect 2964 13132 3016 13184
rect 4804 13132 4856 13184
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 6000 13132 6052 13184
rect 6828 13132 6880 13184
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 8668 13132 8720 13184
rect 9496 13175 9548 13184
rect 9496 13141 9505 13175
rect 9505 13141 9539 13175
rect 9539 13141 9548 13175
rect 9496 13132 9548 13141
rect 10048 13175 10100 13184
rect 10048 13141 10057 13175
rect 10057 13141 10091 13175
rect 10091 13141 10100 13175
rect 10048 13132 10100 13141
rect 10784 13175 10836 13184
rect 10784 13141 10793 13175
rect 10793 13141 10827 13175
rect 10827 13141 10836 13175
rect 10784 13132 10836 13141
rect 11612 13132 11664 13184
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 16488 13175 16540 13184
rect 16488 13141 16497 13175
rect 16497 13141 16531 13175
rect 16531 13141 16540 13175
rect 16488 13132 16540 13141
rect 3696 13030 3748 13082
rect 3760 13030 3812 13082
rect 3824 13030 3876 13082
rect 3888 13030 3940 13082
rect 9124 13030 9176 13082
rect 9188 13030 9240 13082
rect 9252 13030 9304 13082
rect 9316 13030 9368 13082
rect 14552 13030 14604 13082
rect 14616 13030 14668 13082
rect 14680 13030 14732 13082
rect 14744 13030 14796 13082
rect 4620 12928 4672 12980
rect 5172 12928 5224 12980
rect 7840 12971 7892 12980
rect 7840 12937 7849 12971
rect 7849 12937 7883 12971
rect 7883 12937 7892 12971
rect 7840 12928 7892 12937
rect 8668 12971 8720 12980
rect 8668 12937 8677 12971
rect 8677 12937 8711 12971
rect 8711 12937 8720 12971
rect 8668 12928 8720 12937
rect 10140 12928 10192 12980
rect 16396 12971 16448 12980
rect 16396 12937 16405 12971
rect 16405 12937 16439 12971
rect 16439 12937 16448 12971
rect 16396 12928 16448 12937
rect 1492 12835 1544 12844
rect 1492 12801 1501 12835
rect 1501 12801 1535 12835
rect 1535 12801 1544 12835
rect 1492 12792 1544 12801
rect 4528 12860 4580 12912
rect 4988 12860 5040 12912
rect 2872 12792 2924 12844
rect 2780 12724 2832 12776
rect 3056 12656 3108 12708
rect 4160 12724 4212 12776
rect 5264 12767 5316 12776
rect 5264 12733 5273 12767
rect 5273 12733 5307 12767
rect 5307 12733 5316 12767
rect 5264 12724 5316 12733
rect 5540 12724 5592 12776
rect 6000 12767 6052 12776
rect 6000 12733 6009 12767
rect 6009 12733 6043 12767
rect 6043 12733 6052 12767
rect 6000 12724 6052 12733
rect 7288 12656 7340 12708
rect 7932 12656 7984 12708
rect 8576 12724 8628 12776
rect 9772 12792 9824 12844
rect 10692 12792 10744 12844
rect 16580 12792 16632 12844
rect 9404 12767 9456 12776
rect 9404 12733 9413 12767
rect 9413 12733 9447 12767
rect 9447 12733 9456 12767
rect 9404 12724 9456 12733
rect 11336 12724 11388 12776
rect 8484 12656 8536 12708
rect 8668 12656 8720 12708
rect 9680 12699 9732 12708
rect 9680 12665 9689 12699
rect 9689 12665 9723 12699
rect 9723 12665 9732 12699
rect 9680 12656 9732 12665
rect 10416 12656 10468 12708
rect 13636 12656 13688 12708
rect 13912 12699 13964 12708
rect 13912 12665 13921 12699
rect 13921 12665 13955 12699
rect 13955 12665 13964 12699
rect 13912 12656 13964 12665
rect 1860 12631 1912 12640
rect 1860 12597 1869 12631
rect 1869 12597 1903 12631
rect 1903 12597 1912 12631
rect 1860 12588 1912 12597
rect 4068 12631 4120 12640
rect 4068 12597 4077 12631
rect 4077 12597 4111 12631
rect 4111 12597 4120 12631
rect 4068 12588 4120 12597
rect 5264 12588 5316 12640
rect 5816 12631 5868 12640
rect 5816 12597 5825 12631
rect 5825 12597 5859 12631
rect 5859 12597 5868 12631
rect 5816 12588 5868 12597
rect 8024 12588 8076 12640
rect 11428 12588 11480 12640
rect 16028 12724 16080 12776
rect 14924 12656 14976 12708
rect 6410 12486 6462 12538
rect 6474 12486 6526 12538
rect 6538 12486 6590 12538
rect 6602 12486 6654 12538
rect 11838 12486 11890 12538
rect 11902 12486 11954 12538
rect 11966 12486 12018 12538
rect 12030 12486 12082 12538
rect 1400 12427 1452 12436
rect 1400 12393 1409 12427
rect 1409 12393 1443 12427
rect 1443 12393 1452 12427
rect 1400 12384 1452 12393
rect 5540 12384 5592 12436
rect 9588 12384 9640 12436
rect 11704 12427 11756 12436
rect 3056 12359 3108 12368
rect 1860 12248 1912 12300
rect 3056 12325 3065 12359
rect 3065 12325 3099 12359
rect 3099 12325 3108 12359
rect 3056 12316 3108 12325
rect 4804 12359 4856 12368
rect 4804 12325 4813 12359
rect 4813 12325 4847 12359
rect 4847 12325 4856 12359
rect 4804 12316 4856 12325
rect 6920 12316 6972 12368
rect 7748 12316 7800 12368
rect 9956 12316 10008 12368
rect 11704 12393 11713 12427
rect 11713 12393 11747 12427
rect 11747 12393 11756 12427
rect 11704 12384 11756 12393
rect 12440 12384 12492 12436
rect 10600 12316 10652 12368
rect 2136 12248 2188 12300
rect 3516 12248 3568 12300
rect 5908 12248 5960 12300
rect 9496 12291 9548 12300
rect 9496 12257 9505 12291
rect 9505 12257 9539 12291
rect 9539 12257 9548 12291
rect 9496 12248 9548 12257
rect 2228 12180 2280 12232
rect 2964 12180 3016 12232
rect 5540 12180 5592 12232
rect 5816 12180 5868 12232
rect 9864 12291 9916 12300
rect 9864 12257 9873 12291
rect 9873 12257 9907 12291
rect 9907 12257 9916 12291
rect 9864 12248 9916 12257
rect 10140 12180 10192 12232
rect 9680 12112 9732 12164
rect 11612 12248 11664 12300
rect 12348 12248 12400 12300
rect 12900 12384 12952 12436
rect 13636 12427 13688 12436
rect 13636 12393 13645 12427
rect 13645 12393 13679 12427
rect 13679 12393 13688 12427
rect 13636 12384 13688 12393
rect 13912 12384 13964 12436
rect 15200 12316 15252 12368
rect 16396 12384 16448 12436
rect 16580 12427 16632 12436
rect 16580 12393 16589 12427
rect 16589 12393 16623 12427
rect 16623 12393 16632 12427
rect 16580 12384 16632 12393
rect 16212 12359 16264 12368
rect 16212 12325 16221 12359
rect 16221 12325 16255 12359
rect 16255 12325 16264 12359
rect 16212 12316 16264 12325
rect 15936 12248 15988 12300
rect 16488 12248 16540 12300
rect 3516 12044 3568 12096
rect 4344 12044 4396 12096
rect 9864 12044 9916 12096
rect 12072 12044 12124 12096
rect 13360 12044 13412 12096
rect 13820 12044 13872 12096
rect 3696 11942 3748 11994
rect 3760 11942 3812 11994
rect 3824 11942 3876 11994
rect 3888 11942 3940 11994
rect 9124 11942 9176 11994
rect 9188 11942 9240 11994
rect 9252 11942 9304 11994
rect 9316 11942 9368 11994
rect 14552 11942 14604 11994
rect 14616 11942 14668 11994
rect 14680 11942 14732 11994
rect 14744 11942 14796 11994
rect 4620 11883 4672 11892
rect 4620 11849 4629 11883
rect 4629 11849 4663 11883
rect 4663 11849 4672 11883
rect 4620 11840 4672 11849
rect 7748 11883 7800 11892
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 10692 11840 10744 11892
rect 12716 11840 12768 11892
rect 2964 11704 3016 11756
rect 4528 11747 4580 11756
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4528 11704 4580 11713
rect 9496 11704 9548 11756
rect 11428 11704 11480 11756
rect 14924 11704 14976 11756
rect 4068 11636 4120 11688
rect 7564 11679 7616 11688
rect 7564 11645 7573 11679
rect 7573 11645 7607 11679
rect 7607 11645 7616 11679
rect 7564 11636 7616 11645
rect 10600 11636 10652 11688
rect 12072 11679 12124 11688
rect 12072 11645 12081 11679
rect 12081 11645 12115 11679
rect 12115 11645 12124 11679
rect 12072 11636 12124 11645
rect 12348 11679 12400 11688
rect 12348 11645 12357 11679
rect 12357 11645 12391 11679
rect 12391 11645 12400 11679
rect 12348 11636 12400 11645
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 16396 11679 16448 11688
rect 12440 11636 12492 11645
rect 16396 11645 16405 11679
rect 16405 11645 16439 11679
rect 16439 11645 16448 11679
rect 16396 11636 16448 11645
rect 2596 11611 2648 11620
rect 2596 11577 2605 11611
rect 2605 11577 2639 11611
rect 2639 11577 2648 11611
rect 2596 11568 2648 11577
rect 12256 11611 12308 11620
rect 12256 11577 12265 11611
rect 12265 11577 12299 11611
rect 12299 11577 12308 11611
rect 12256 11568 12308 11577
rect 13820 11568 13872 11620
rect 15476 11611 15528 11620
rect 15476 11577 15485 11611
rect 15485 11577 15519 11611
rect 15519 11577 15528 11611
rect 15476 11568 15528 11577
rect 2688 11500 2740 11552
rect 4620 11500 4672 11552
rect 5080 11500 5132 11552
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 10692 11500 10744 11552
rect 14004 11543 14056 11552
rect 14004 11509 14013 11543
rect 14013 11509 14047 11543
rect 14047 11509 14056 11543
rect 14004 11500 14056 11509
rect 16212 11543 16264 11552
rect 16212 11509 16221 11543
rect 16221 11509 16255 11543
rect 16255 11509 16264 11543
rect 16212 11500 16264 11509
rect 6410 11398 6462 11450
rect 6474 11398 6526 11450
rect 6538 11398 6590 11450
rect 6602 11398 6654 11450
rect 11838 11398 11890 11450
rect 11902 11398 11954 11450
rect 11966 11398 12018 11450
rect 12030 11398 12082 11450
rect 2136 11339 2188 11348
rect 2136 11305 2145 11339
rect 2145 11305 2179 11339
rect 2179 11305 2188 11339
rect 2136 11296 2188 11305
rect 2412 11296 2464 11348
rect 1768 11203 1820 11212
rect 1768 11169 1777 11203
rect 1777 11169 1811 11203
rect 1811 11169 1820 11203
rect 1768 11160 1820 11169
rect 2320 11203 2372 11212
rect 2320 11169 2326 11203
rect 2326 11169 2360 11203
rect 2360 11169 2372 11203
rect 2320 11160 2372 11169
rect 2688 11160 2740 11212
rect 5632 11296 5684 11348
rect 7472 11296 7524 11348
rect 12164 11296 12216 11348
rect 13820 11339 13872 11348
rect 13820 11305 13829 11339
rect 13829 11305 13863 11339
rect 13863 11305 13872 11339
rect 13820 11296 13872 11305
rect 16488 11296 16540 11348
rect 5080 11228 5132 11280
rect 5816 11228 5868 11280
rect 9588 11228 9640 11280
rect 11336 11228 11388 11280
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 12256 11203 12308 11212
rect 12256 11169 12268 11203
rect 12268 11169 12302 11203
rect 12302 11169 12308 11203
rect 12256 11160 12308 11169
rect 13360 11160 13412 11212
rect 15200 11228 15252 11280
rect 16212 11228 16264 11280
rect 14924 11203 14976 11212
rect 14924 11169 14933 11203
rect 14933 11169 14967 11203
rect 14967 11169 14976 11203
rect 14924 11160 14976 11169
rect 4068 11092 4120 11144
rect 5540 11092 5592 11144
rect 7380 11092 7432 11144
rect 10600 11092 10652 11144
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 11428 11092 11480 11144
rect 11704 11092 11756 11144
rect 7472 11067 7524 11076
rect 7472 11033 7481 11067
rect 7481 11033 7515 11067
rect 7515 11033 7524 11067
rect 7472 11024 7524 11033
rect 8392 11067 8444 11076
rect 8392 11033 8401 11067
rect 8401 11033 8435 11067
rect 8435 11033 8444 11067
rect 8392 11024 8444 11033
rect 13084 11067 13136 11076
rect 13084 11033 13093 11067
rect 13093 11033 13127 11067
rect 13127 11033 13136 11067
rect 13084 11024 13136 11033
rect 2412 10956 2464 11008
rect 7012 10956 7064 11008
rect 7104 10956 7156 11008
rect 7564 10956 7616 11008
rect 10876 10956 10928 11008
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 15200 10999 15252 11008
rect 12440 10956 12492 10965
rect 15200 10965 15230 10999
rect 15230 10965 15252 10999
rect 15200 10956 15252 10965
rect 3696 10854 3748 10906
rect 3760 10854 3812 10906
rect 3824 10854 3876 10906
rect 3888 10854 3940 10906
rect 9124 10854 9176 10906
rect 9188 10854 9240 10906
rect 9252 10854 9304 10906
rect 9316 10854 9368 10906
rect 14552 10854 14604 10906
rect 14616 10854 14668 10906
rect 14680 10854 14732 10906
rect 14744 10854 14796 10906
rect 2596 10795 2648 10804
rect 2596 10761 2605 10795
rect 2605 10761 2639 10795
rect 2639 10761 2648 10795
rect 2596 10752 2648 10761
rect 4068 10752 4120 10804
rect 5264 10752 5316 10804
rect 10048 10752 10100 10804
rect 11060 10752 11112 10804
rect 11336 10795 11388 10804
rect 11336 10761 11345 10795
rect 11345 10761 11379 10795
rect 11379 10761 11388 10795
rect 11336 10752 11388 10761
rect 15476 10752 15528 10804
rect 13636 10684 13688 10736
rect 2136 10548 2188 10600
rect 2228 10591 2280 10600
rect 2228 10557 2237 10591
rect 2237 10557 2271 10591
rect 2271 10557 2280 10591
rect 2412 10591 2464 10600
rect 2228 10548 2280 10557
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 3240 10591 3292 10600
rect 3240 10557 3249 10591
rect 3249 10557 3283 10591
rect 3283 10557 3292 10591
rect 3240 10548 3292 10557
rect 5080 10548 5132 10600
rect 9496 10548 9548 10600
rect 9680 10591 9732 10600
rect 11428 10616 11480 10668
rect 12440 10616 12492 10668
rect 9680 10557 9722 10591
rect 9722 10557 9732 10591
rect 9680 10548 9732 10557
rect 10692 10591 10744 10600
rect 2320 10523 2372 10532
rect 2320 10489 2329 10523
rect 2329 10489 2363 10523
rect 2363 10489 2372 10523
rect 2320 10480 2372 10489
rect 8392 10480 8444 10532
rect 8852 10523 8904 10532
rect 8852 10489 8861 10523
rect 8861 10489 8895 10523
rect 8895 10489 8904 10523
rect 8852 10480 8904 10489
rect 3056 10455 3108 10464
rect 3056 10421 3065 10455
rect 3065 10421 3099 10455
rect 3099 10421 3108 10455
rect 3056 10412 3108 10421
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 10048 10480 10100 10532
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 10692 10548 10744 10557
rect 10784 10548 10836 10600
rect 10600 10523 10652 10532
rect 10600 10489 10609 10523
rect 10609 10489 10643 10523
rect 10643 10489 10652 10523
rect 10600 10480 10652 10489
rect 13084 10480 13136 10532
rect 14004 10548 14056 10600
rect 14924 10455 14976 10464
rect 14924 10421 14933 10455
rect 14933 10421 14967 10455
rect 14967 10421 14976 10455
rect 14924 10412 14976 10421
rect 6410 10310 6462 10362
rect 6474 10310 6526 10362
rect 6538 10310 6590 10362
rect 6602 10310 6654 10362
rect 11838 10310 11890 10362
rect 11902 10310 11954 10362
rect 11966 10310 12018 10362
rect 12030 10310 12082 10362
rect 3332 10208 3384 10260
rect 5080 10208 5132 10260
rect 5816 10251 5868 10260
rect 5816 10217 5825 10251
rect 5825 10217 5859 10251
rect 5859 10217 5868 10251
rect 5816 10208 5868 10217
rect 6920 10208 6972 10260
rect 7012 10251 7064 10260
rect 7012 10217 7021 10251
rect 7021 10217 7055 10251
rect 7055 10217 7064 10251
rect 7012 10208 7064 10217
rect 1400 10140 1452 10192
rect 3056 10140 3108 10192
rect 7104 10140 7156 10192
rect 7472 10208 7524 10260
rect 7380 10140 7432 10192
rect 2964 10004 3016 10056
rect 8116 10115 8168 10124
rect 8116 10081 8125 10115
rect 8125 10081 8159 10115
rect 8159 10081 8168 10115
rect 8116 10072 8168 10081
rect 8852 10208 8904 10260
rect 11704 10251 11756 10260
rect 11704 10217 11713 10251
rect 11713 10217 11747 10251
rect 11747 10217 11756 10251
rect 11704 10208 11756 10217
rect 8944 10072 8996 10124
rect 11152 10072 11204 10124
rect 12808 10072 12860 10124
rect 13176 10115 13228 10124
rect 13176 10081 13182 10115
rect 13182 10081 13216 10115
rect 13216 10081 13228 10115
rect 15752 10140 15804 10192
rect 13176 10072 13228 10081
rect 14924 10072 14976 10124
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 15568 10115 15620 10124
rect 15568 10081 15577 10115
rect 15577 10081 15611 10115
rect 15611 10081 15620 10115
rect 15844 10115 15896 10124
rect 15568 10072 15620 10081
rect 15844 10081 15853 10115
rect 15853 10081 15887 10115
rect 15887 10081 15896 10115
rect 15844 10072 15896 10081
rect 16396 10072 16448 10124
rect 13636 10047 13688 10056
rect 13636 10013 13645 10047
rect 13645 10013 13679 10047
rect 13679 10013 13688 10047
rect 13636 10004 13688 10013
rect 8484 9936 8536 9988
rect 9496 9936 9548 9988
rect 13268 9868 13320 9920
rect 15292 9911 15344 9920
rect 15292 9877 15301 9911
rect 15301 9877 15335 9911
rect 15335 9877 15344 9911
rect 15292 9868 15344 9877
rect 16304 9911 16356 9920
rect 16304 9877 16313 9911
rect 16313 9877 16347 9911
rect 16347 9877 16356 9911
rect 16304 9868 16356 9877
rect 3696 9766 3748 9818
rect 3760 9766 3812 9818
rect 3824 9766 3876 9818
rect 3888 9766 3940 9818
rect 9124 9766 9176 9818
rect 9188 9766 9240 9818
rect 9252 9766 9304 9818
rect 9316 9766 9368 9818
rect 14552 9766 14604 9818
rect 14616 9766 14668 9818
rect 14680 9766 14732 9818
rect 14744 9766 14796 9818
rect 15844 9707 15896 9716
rect 3240 9460 3292 9512
rect 4712 9460 4764 9512
rect 5264 9503 5316 9512
rect 5264 9469 5273 9503
rect 5273 9469 5307 9503
rect 5307 9469 5316 9503
rect 5264 9460 5316 9469
rect 6276 9596 6328 9648
rect 7196 9596 7248 9648
rect 15844 9673 15853 9707
rect 15853 9673 15887 9707
rect 15887 9673 15896 9707
rect 15844 9664 15896 9673
rect 7104 9460 7156 9512
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 10600 9596 10652 9648
rect 9956 9571 10008 9580
rect 9956 9537 9965 9571
rect 9965 9537 9999 9571
rect 9999 9537 10008 9571
rect 12348 9596 12400 9648
rect 9956 9528 10008 9537
rect 10600 9503 10652 9512
rect 10600 9469 10606 9503
rect 10606 9469 10640 9503
rect 10640 9469 10652 9503
rect 10600 9460 10652 9469
rect 3516 9324 3568 9376
rect 4712 9324 4764 9376
rect 10508 9392 10560 9444
rect 6828 9367 6880 9376
rect 6828 9333 6837 9367
rect 6837 9333 6871 9367
rect 6871 9333 6880 9367
rect 6828 9324 6880 9333
rect 7196 9324 7248 9376
rect 10416 9367 10468 9376
rect 10416 9333 10425 9367
rect 10425 9333 10459 9367
rect 10459 9333 10468 9367
rect 10416 9324 10468 9333
rect 13268 9571 13320 9580
rect 12440 9460 12492 9512
rect 12164 9324 12216 9376
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 13820 9392 13872 9444
rect 14924 9324 14976 9376
rect 15476 9528 15528 9580
rect 15568 9460 15620 9512
rect 15936 9460 15988 9512
rect 6410 9222 6462 9274
rect 6474 9222 6526 9274
rect 6538 9222 6590 9274
rect 6602 9222 6654 9274
rect 11838 9222 11890 9274
rect 11902 9222 11954 9274
rect 11966 9222 12018 9274
rect 12030 9222 12082 9274
rect 1400 9163 1452 9172
rect 1400 9129 1409 9163
rect 1409 9129 1443 9163
rect 1443 9129 1452 9163
rect 1400 9120 1452 9129
rect 2688 9163 2740 9172
rect 1860 8984 1912 9036
rect 2688 9129 2697 9163
rect 2697 9129 2731 9163
rect 2731 9129 2740 9163
rect 2688 9120 2740 9129
rect 7104 9120 7156 9172
rect 7472 9120 7524 9172
rect 4712 9052 4764 9104
rect 10600 9120 10652 9172
rect 13176 9163 13228 9172
rect 13176 9129 13185 9163
rect 13185 9129 13219 9163
rect 13219 9129 13228 9163
rect 13176 9120 13228 9129
rect 13820 9163 13872 9172
rect 13820 9129 13829 9163
rect 13829 9129 13863 9163
rect 13863 9129 13872 9163
rect 13820 9120 13872 9129
rect 15936 9120 15988 9172
rect 12164 9052 12216 9104
rect 15292 9052 15344 9104
rect 2596 8984 2648 9036
rect 7840 8984 7892 9036
rect 9772 9027 9824 9036
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 2320 8780 2372 8832
rect 2688 8780 2740 8832
rect 6276 8916 6328 8968
rect 7380 8916 7432 8968
rect 9772 8993 9781 9027
rect 9781 8993 9815 9027
rect 9815 8993 9824 9027
rect 9772 8984 9824 8993
rect 9956 9027 10008 9036
rect 9956 8993 9965 9027
rect 9965 8993 9999 9027
rect 9999 8993 10008 9027
rect 9956 8984 10008 8993
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 13360 8984 13412 9036
rect 14924 9027 14976 9036
rect 14924 8993 14933 9027
rect 14933 8993 14967 9027
rect 14967 8993 14976 9027
rect 14924 8984 14976 8993
rect 16304 8984 16356 9036
rect 10416 8916 10468 8968
rect 10600 8959 10652 8968
rect 10600 8925 10609 8959
rect 10609 8925 10643 8959
rect 10643 8925 10652 8959
rect 10600 8916 10652 8925
rect 12808 8959 12860 8968
rect 12808 8925 12817 8959
rect 12817 8925 12851 8959
rect 12851 8925 12860 8959
rect 12808 8916 12860 8925
rect 13728 8916 13780 8968
rect 8024 8780 8076 8832
rect 3696 8678 3748 8730
rect 3760 8678 3812 8730
rect 3824 8678 3876 8730
rect 3888 8678 3940 8730
rect 9124 8678 9176 8730
rect 9188 8678 9240 8730
rect 9252 8678 9304 8730
rect 9316 8678 9368 8730
rect 14552 8678 14604 8730
rect 14616 8678 14668 8730
rect 14680 8678 14732 8730
rect 14744 8678 14796 8730
rect 2596 8619 2648 8628
rect 2596 8585 2605 8619
rect 2605 8585 2639 8619
rect 2639 8585 2648 8619
rect 2596 8576 2648 8585
rect 4712 8508 4764 8560
rect 6276 8576 6328 8628
rect 7380 8619 7432 8628
rect 7380 8585 7389 8619
rect 7389 8585 7423 8619
rect 7423 8585 7432 8619
rect 7380 8576 7432 8585
rect 8116 8576 8168 8628
rect 9680 8576 9732 8628
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 10508 8576 10560 8628
rect 12808 8576 12860 8628
rect 5448 8508 5500 8560
rect 15200 8576 15252 8628
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 3516 8304 3568 8356
rect 4068 8347 4120 8356
rect 4068 8313 4077 8347
rect 4077 8313 4111 8347
rect 4111 8313 4120 8347
rect 4068 8304 4120 8313
rect 4344 8304 4396 8356
rect 4712 8304 4764 8356
rect 7288 8440 7340 8492
rect 5448 8372 5500 8424
rect 5816 8372 5868 8424
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 7104 8415 7156 8424
rect 7104 8381 7113 8415
rect 7113 8381 7147 8415
rect 7147 8381 7156 8415
rect 7104 8372 7156 8381
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 2044 8236 2096 8288
rect 2504 8236 2556 8288
rect 5356 8304 5408 8356
rect 15476 8508 15528 8560
rect 8760 8440 8812 8492
rect 8576 8304 8628 8356
rect 9772 8372 9824 8424
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 13544 8440 13596 8492
rect 14924 8440 14976 8492
rect 12164 8372 12216 8424
rect 15568 8372 15620 8424
rect 10416 8304 10468 8356
rect 13820 8304 13872 8356
rect 15844 8576 15896 8628
rect 15752 8508 15804 8560
rect 16396 8415 16448 8424
rect 16396 8381 16405 8415
rect 16405 8381 16439 8415
rect 16439 8381 16448 8415
rect 16396 8372 16448 8381
rect 6276 8279 6328 8288
rect 6276 8245 6285 8279
rect 6285 8245 6319 8279
rect 6319 8245 6328 8279
rect 6276 8236 6328 8245
rect 6736 8236 6788 8288
rect 9956 8236 10008 8288
rect 10600 8236 10652 8288
rect 12348 8236 12400 8288
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 15844 8236 15896 8288
rect 6410 8134 6462 8186
rect 6474 8134 6526 8186
rect 6538 8134 6590 8186
rect 6602 8134 6654 8186
rect 11838 8134 11890 8186
rect 11902 8134 11954 8186
rect 11966 8134 12018 8186
rect 12030 8134 12082 8186
rect 1676 8032 1728 8084
rect 4068 8032 4120 8084
rect 5356 8032 5408 8084
rect 2596 8007 2648 8016
rect 2596 7973 2605 8007
rect 2605 7973 2639 8007
rect 2639 7973 2648 8007
rect 2596 7964 2648 7973
rect 1952 7939 2004 7948
rect 1952 7905 1961 7939
rect 1961 7905 1995 7939
rect 1995 7905 2004 7939
rect 1952 7896 2004 7905
rect 2320 7939 2372 7948
rect 2320 7905 2329 7939
rect 2329 7905 2363 7939
rect 2363 7905 2372 7939
rect 2320 7896 2372 7905
rect 2504 7939 2556 7948
rect 2504 7905 2513 7939
rect 2513 7905 2547 7939
rect 2547 7905 2556 7939
rect 2504 7896 2556 7905
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 4620 7964 4672 8016
rect 7840 7964 7892 8016
rect 11060 8032 11112 8084
rect 8760 7964 8812 8016
rect 9956 7964 10008 8016
rect 10784 7964 10836 8016
rect 12532 8032 12584 8084
rect 13820 8075 13872 8084
rect 13820 8041 13829 8075
rect 13829 8041 13863 8075
rect 13863 8041 13872 8075
rect 13820 8032 13872 8041
rect 14924 8075 14976 8084
rect 14924 8041 14933 8075
rect 14933 8041 14967 8075
rect 14967 8041 14976 8075
rect 14924 8032 14976 8041
rect 15660 8032 15712 8084
rect 12440 7964 12492 8016
rect 13176 7964 13228 8016
rect 4528 7939 4580 7948
rect 4528 7905 4537 7939
rect 4537 7905 4571 7939
rect 4571 7905 4580 7939
rect 4528 7896 4580 7905
rect 4712 7896 4764 7948
rect 9496 7939 9548 7948
rect 9496 7905 9505 7939
rect 9505 7905 9539 7939
rect 9539 7905 9548 7939
rect 9496 7896 9548 7905
rect 13728 7964 13780 8016
rect 5448 7828 5500 7880
rect 10600 7828 10652 7880
rect 12808 7828 12860 7880
rect 13084 7828 13136 7880
rect 12256 7760 12308 7812
rect 15292 7896 15344 7948
rect 16672 7939 16724 7948
rect 16672 7905 16681 7939
rect 16681 7905 16715 7939
rect 16715 7905 16724 7939
rect 16672 7896 16724 7905
rect 15476 7760 15528 7812
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 9680 7735 9732 7744
rect 9680 7701 9689 7735
rect 9689 7701 9723 7735
rect 9723 7701 9732 7735
rect 9680 7692 9732 7701
rect 10416 7692 10468 7744
rect 12164 7692 12216 7744
rect 12532 7735 12584 7744
rect 12532 7701 12541 7735
rect 12541 7701 12575 7735
rect 12575 7701 12584 7735
rect 12532 7692 12584 7701
rect 13360 7692 13412 7744
rect 3696 7590 3748 7642
rect 3760 7590 3812 7642
rect 3824 7590 3876 7642
rect 3888 7590 3940 7642
rect 9124 7590 9176 7642
rect 9188 7590 9240 7642
rect 9252 7590 9304 7642
rect 9316 7590 9368 7642
rect 14552 7590 14604 7642
rect 14616 7590 14668 7642
rect 14680 7590 14732 7642
rect 14744 7590 14796 7642
rect 3516 7488 3568 7540
rect 4068 7488 4120 7540
rect 5448 7488 5500 7540
rect 10508 7531 10560 7540
rect 1676 7148 1728 7200
rect 4252 7352 4304 7404
rect 3148 7284 3200 7336
rect 4068 7284 4120 7336
rect 5816 7420 5868 7472
rect 7656 7420 7708 7472
rect 8484 7420 8536 7472
rect 5724 7352 5776 7404
rect 7012 7327 7064 7336
rect 7012 7293 7021 7327
rect 7021 7293 7055 7327
rect 7055 7293 7064 7327
rect 7012 7284 7064 7293
rect 8208 7327 8260 7336
rect 8208 7293 8220 7327
rect 8220 7293 8254 7327
rect 8254 7293 8260 7327
rect 8208 7284 8260 7293
rect 9680 7352 9732 7404
rect 10508 7497 10517 7531
rect 10517 7497 10551 7531
rect 10551 7497 10560 7531
rect 10508 7488 10560 7497
rect 10784 7488 10836 7540
rect 12072 7395 12124 7404
rect 12072 7361 12081 7395
rect 12081 7361 12115 7395
rect 12115 7361 12124 7395
rect 12072 7352 12124 7361
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 10324 7327 10376 7336
rect 10324 7293 10333 7327
rect 10333 7293 10367 7327
rect 10367 7293 10376 7327
rect 10324 7284 10376 7293
rect 11060 7284 11112 7336
rect 16212 7352 16264 7404
rect 12348 7284 12400 7336
rect 15844 7327 15896 7336
rect 15844 7293 15853 7327
rect 15853 7293 15887 7327
rect 15887 7293 15896 7327
rect 15844 7284 15896 7293
rect 15936 7327 15988 7336
rect 15936 7293 15945 7327
rect 15945 7293 15979 7327
rect 15979 7293 15988 7327
rect 15936 7284 15988 7293
rect 13268 7259 13320 7268
rect 13268 7225 13277 7259
rect 13277 7225 13311 7259
rect 13311 7225 13320 7259
rect 13268 7216 13320 7225
rect 13820 7216 13872 7268
rect 3516 7148 3568 7200
rect 4252 7191 4304 7200
rect 4252 7157 4261 7191
rect 4261 7157 4295 7191
rect 4295 7157 4304 7191
rect 4252 7148 4304 7157
rect 4804 7148 4856 7200
rect 5448 7191 5500 7200
rect 5448 7157 5457 7191
rect 5457 7157 5491 7191
rect 5491 7157 5500 7191
rect 5448 7148 5500 7157
rect 6092 7148 6144 7200
rect 7656 7148 7708 7200
rect 8484 7148 8536 7200
rect 9496 7191 9548 7200
rect 9496 7157 9505 7191
rect 9505 7157 9539 7191
rect 9539 7157 9548 7191
rect 9496 7148 9548 7157
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 15016 7148 15068 7200
rect 6410 7046 6462 7098
rect 6474 7046 6526 7098
rect 6538 7046 6590 7098
rect 6602 7046 6654 7098
rect 11838 7046 11890 7098
rect 11902 7046 11954 7098
rect 11966 7046 12018 7098
rect 12030 7046 12082 7098
rect 7012 6944 7064 6996
rect 1676 6919 1728 6928
rect 1676 6885 1685 6919
rect 1685 6885 1719 6919
rect 1719 6885 1728 6919
rect 1676 6876 1728 6885
rect 2412 6876 2464 6928
rect 4804 6919 4856 6928
rect 4804 6885 4813 6919
rect 4813 6885 4847 6919
rect 4847 6885 4856 6919
rect 4804 6876 4856 6885
rect 6092 6876 6144 6928
rect 6736 6851 6788 6860
rect 6736 6817 6745 6851
rect 6745 6817 6779 6851
rect 6779 6817 6788 6851
rect 6736 6808 6788 6817
rect 2044 6740 2096 6792
rect 2320 6740 2372 6792
rect 4896 6740 4948 6792
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 8208 6740 8260 6792
rect 12164 6944 12216 6996
rect 13268 6944 13320 6996
rect 10416 6808 10468 6860
rect 12440 6808 12492 6860
rect 12164 6740 12216 6792
rect 13084 6808 13136 6860
rect 13360 6851 13412 6860
rect 13360 6817 13369 6851
rect 13369 6817 13403 6851
rect 13403 6817 13412 6851
rect 13360 6808 13412 6817
rect 14924 6808 14976 6860
rect 10600 6672 10652 6724
rect 13544 6715 13596 6724
rect 7656 6604 7708 6656
rect 9772 6604 9824 6656
rect 12256 6604 12308 6656
rect 13544 6681 13553 6715
rect 13553 6681 13587 6715
rect 13587 6681 13596 6715
rect 13544 6672 13596 6681
rect 14372 6672 14424 6724
rect 15384 6851 15436 6860
rect 15384 6817 15393 6851
rect 15393 6817 15427 6851
rect 15427 6817 15436 6851
rect 15384 6808 15436 6817
rect 15568 6808 15620 6860
rect 16120 6808 16172 6860
rect 15660 6740 15712 6792
rect 15936 6740 15988 6792
rect 15108 6604 15160 6656
rect 15200 6604 15252 6656
rect 3696 6502 3748 6554
rect 3760 6502 3812 6554
rect 3824 6502 3876 6554
rect 3888 6502 3940 6554
rect 9124 6502 9176 6554
rect 9188 6502 9240 6554
rect 9252 6502 9304 6554
rect 9316 6502 9368 6554
rect 14552 6502 14604 6554
rect 14616 6502 14668 6554
rect 14680 6502 14732 6554
rect 14744 6502 14796 6554
rect 2412 6443 2464 6452
rect 2412 6409 2421 6443
rect 2421 6409 2455 6443
rect 2455 6409 2464 6443
rect 2412 6400 2464 6409
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 7012 6400 7064 6452
rect 4252 6264 4304 6316
rect 11152 6400 11204 6452
rect 13820 6400 13872 6452
rect 14924 6443 14976 6452
rect 2780 6196 2832 6248
rect 4896 6239 4948 6248
rect 4896 6205 4905 6239
rect 4905 6205 4939 6239
rect 4939 6205 4948 6239
rect 4896 6196 4948 6205
rect 5172 6196 5224 6248
rect 4160 6128 4212 6180
rect 1584 6060 1636 6112
rect 9404 6264 9456 6316
rect 5632 6196 5684 6248
rect 7104 6239 7156 6248
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 7656 6196 7708 6248
rect 8208 6239 8260 6248
rect 8208 6205 8217 6239
rect 8217 6205 8251 6239
rect 8251 6205 8260 6239
rect 8484 6239 8536 6248
rect 8208 6196 8260 6205
rect 8484 6205 8493 6239
rect 8493 6205 8527 6239
rect 8527 6205 8536 6239
rect 8484 6196 8536 6205
rect 8852 6128 8904 6180
rect 5724 6103 5776 6112
rect 5724 6069 5733 6103
rect 5733 6069 5767 6103
rect 5767 6069 5776 6103
rect 5724 6060 5776 6069
rect 6920 6103 6972 6112
rect 6920 6069 6929 6103
rect 6929 6069 6963 6103
rect 6963 6069 6972 6103
rect 6920 6060 6972 6069
rect 12256 6196 12308 6248
rect 13176 6239 13228 6248
rect 13176 6205 13185 6239
rect 13185 6205 13219 6239
rect 13219 6205 13228 6239
rect 13176 6196 13228 6205
rect 14372 6239 14424 6248
rect 14372 6205 14382 6239
rect 14382 6205 14424 6239
rect 14372 6196 14424 6205
rect 9772 6128 9824 6180
rect 14924 6409 14933 6443
rect 14933 6409 14967 6443
rect 14967 6409 14976 6443
rect 14924 6400 14976 6409
rect 15016 6400 15068 6452
rect 15568 6400 15620 6452
rect 16212 6443 16264 6452
rect 16212 6409 16221 6443
rect 16221 6409 16255 6443
rect 16255 6409 16264 6443
rect 16212 6400 16264 6409
rect 15384 6196 15436 6248
rect 15568 6239 15620 6248
rect 15568 6205 15577 6239
rect 15577 6205 15611 6239
rect 15611 6205 15620 6239
rect 15568 6196 15620 6205
rect 16396 6239 16448 6248
rect 16396 6205 16405 6239
rect 16405 6205 16439 6239
rect 16439 6205 16448 6239
rect 16396 6196 16448 6205
rect 10232 6060 10284 6112
rect 11520 6060 11572 6112
rect 12164 6060 12216 6112
rect 14096 6060 14148 6112
rect 14372 6060 14424 6112
rect 15016 6060 15068 6112
rect 6410 5958 6462 6010
rect 6474 5958 6526 6010
rect 6538 5958 6590 6010
rect 6602 5958 6654 6010
rect 11838 5958 11890 6010
rect 11902 5958 11954 6010
rect 11966 5958 12018 6010
rect 12030 5958 12082 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 4160 5856 4212 5908
rect 4896 5856 4948 5908
rect 6920 5788 6972 5840
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 4068 5720 4120 5772
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 7380 5695 7432 5704
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 10324 5856 10376 5908
rect 11520 5899 11572 5908
rect 8668 5788 8720 5840
rect 11520 5865 11529 5899
rect 11529 5865 11563 5899
rect 11563 5865 11572 5899
rect 11520 5856 11572 5865
rect 15292 5856 15344 5908
rect 15568 5856 15620 5908
rect 15200 5831 15252 5840
rect 10600 5720 10652 5772
rect 10692 5720 10744 5772
rect 7748 5652 7800 5704
rect 9772 5652 9824 5704
rect 15200 5797 15209 5831
rect 15209 5797 15243 5831
rect 15243 5797 15252 5831
rect 15200 5788 15252 5797
rect 16212 5788 16264 5840
rect 12716 5763 12768 5772
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 12808 5763 12860 5772
rect 12808 5729 12817 5763
rect 12817 5729 12851 5763
rect 12851 5729 12860 5763
rect 12808 5720 12860 5729
rect 11060 5584 11112 5636
rect 5908 5559 5960 5568
rect 5908 5525 5917 5559
rect 5917 5525 5951 5559
rect 5951 5525 5960 5559
rect 5908 5516 5960 5525
rect 8208 5559 8260 5568
rect 8208 5525 8217 5559
rect 8217 5525 8251 5559
rect 8251 5525 8260 5559
rect 8208 5516 8260 5525
rect 10600 5516 10652 5568
rect 12440 5559 12492 5568
rect 12440 5525 12449 5559
rect 12449 5525 12483 5559
rect 12483 5525 12492 5559
rect 14096 5652 14148 5704
rect 12440 5516 12492 5525
rect 15936 5516 15988 5568
rect 3696 5414 3748 5466
rect 3760 5414 3812 5466
rect 3824 5414 3876 5466
rect 3888 5414 3940 5466
rect 9124 5414 9176 5466
rect 9188 5414 9240 5466
rect 9252 5414 9304 5466
rect 9316 5414 9368 5466
rect 14552 5414 14604 5466
rect 14616 5414 14668 5466
rect 14680 5414 14732 5466
rect 14744 5414 14796 5466
rect 3516 5312 3568 5364
rect 4528 5312 4580 5364
rect 4804 5312 4856 5364
rect 5448 5312 5500 5364
rect 6092 5312 6144 5364
rect 7380 5312 7432 5364
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 12716 5312 12768 5364
rect 14372 5312 14424 5364
rect 5724 5244 5776 5296
rect 6000 5176 6052 5228
rect 1952 5151 2004 5160
rect 1952 5117 1961 5151
rect 1961 5117 1995 5151
rect 1995 5117 2004 5151
rect 1952 5108 2004 5117
rect 4344 5108 4396 5160
rect 2228 5083 2280 5092
rect 2228 5049 2237 5083
rect 2237 5049 2271 5083
rect 2271 5049 2280 5083
rect 2228 5040 2280 5049
rect 2964 5040 3016 5092
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 10232 5176 10284 5228
rect 11244 5176 11296 5228
rect 12072 5219 12124 5228
rect 12072 5185 12081 5219
rect 12081 5185 12115 5219
rect 12115 5185 12124 5219
rect 12072 5176 12124 5185
rect 12440 5176 12492 5228
rect 14096 5176 14148 5228
rect 5908 5108 5960 5117
rect 6000 4972 6052 5024
rect 6092 4972 6144 5024
rect 7748 5108 7800 5160
rect 8484 5040 8536 5092
rect 9496 5040 9548 5092
rect 12624 5040 12676 5092
rect 13360 5040 13412 5092
rect 15016 5040 15068 5092
rect 9680 5015 9732 5024
rect 9680 4981 9689 5015
rect 9689 4981 9723 5015
rect 9723 4981 9732 5015
rect 9680 4972 9732 4981
rect 10508 5015 10560 5024
rect 10508 4981 10517 5015
rect 10517 4981 10551 5015
rect 10551 4981 10560 5015
rect 10508 4972 10560 4981
rect 11060 4972 11112 5024
rect 16028 5015 16080 5024
rect 16028 4981 16037 5015
rect 16037 4981 16071 5015
rect 16071 4981 16080 5015
rect 16028 4972 16080 4981
rect 6410 4870 6462 4922
rect 6474 4870 6526 4922
rect 6538 4870 6590 4922
rect 6602 4870 6654 4922
rect 11838 4870 11890 4922
rect 11902 4870 11954 4922
rect 11966 4870 12018 4922
rect 12030 4870 12082 4922
rect 2964 4811 3016 4820
rect 2964 4777 2973 4811
rect 2973 4777 3007 4811
rect 3007 4777 3016 4811
rect 2964 4768 3016 4777
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 2780 4632 2832 4641
rect 4068 4632 4120 4684
rect 4896 4768 4948 4820
rect 6000 4811 6052 4820
rect 6000 4777 6009 4811
rect 6009 4777 6043 4811
rect 6043 4777 6052 4811
rect 6000 4768 6052 4777
rect 9496 4811 9548 4820
rect 9496 4777 9505 4811
rect 9505 4777 9539 4811
rect 9539 4777 9548 4811
rect 9496 4768 9548 4777
rect 12808 4811 12860 4820
rect 12808 4777 12817 4811
rect 12817 4777 12851 4811
rect 12851 4777 12860 4811
rect 12808 4768 12860 4777
rect 13360 4768 13412 4820
rect 15016 4768 15068 4820
rect 16212 4811 16264 4820
rect 16212 4777 16221 4811
rect 16221 4777 16255 4811
rect 16255 4777 16264 4811
rect 16212 4768 16264 4777
rect 1952 4564 2004 4616
rect 5632 4632 5684 4684
rect 4528 4607 4580 4616
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 4896 4564 4948 4616
rect 9772 4700 9824 4752
rect 10508 4743 10560 4752
rect 10508 4709 10517 4743
rect 10517 4709 10551 4743
rect 10551 4709 10560 4743
rect 10508 4700 10560 4709
rect 12072 4700 12124 4752
rect 7104 4632 7156 4684
rect 8392 4632 8444 4684
rect 8668 4632 8720 4684
rect 10232 4675 10284 4684
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 4068 4428 4120 4480
rect 8024 4496 8076 4548
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 9772 4564 9824 4616
rect 13360 4632 13412 4684
rect 15200 4632 15252 4684
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 16396 4675 16448 4684
rect 16396 4641 16405 4675
rect 16405 4641 16439 4675
rect 16439 4641 16448 4675
rect 16396 4632 16448 4641
rect 13820 4564 13872 4616
rect 6920 4428 6972 4480
rect 12164 4428 12216 4480
rect 15660 4428 15712 4480
rect 3696 4326 3748 4378
rect 3760 4326 3812 4378
rect 3824 4326 3876 4378
rect 3888 4326 3940 4378
rect 9124 4326 9176 4378
rect 9188 4326 9240 4378
rect 9252 4326 9304 4378
rect 9316 4326 9368 4378
rect 14552 4326 14604 4378
rect 14616 4326 14668 4378
rect 14680 4326 14732 4378
rect 14744 4326 14796 4378
rect 5632 4267 5684 4276
rect 5632 4233 5641 4267
rect 5641 4233 5675 4267
rect 5675 4233 5684 4267
rect 5632 4224 5684 4233
rect 8024 4267 8076 4276
rect 8024 4233 8033 4267
rect 8033 4233 8067 4267
rect 8067 4233 8076 4267
rect 8024 4224 8076 4233
rect 8484 4224 8536 4276
rect 12072 4267 12124 4276
rect 12072 4233 12081 4267
rect 12081 4233 12115 4267
rect 12115 4233 12124 4267
rect 12072 4224 12124 4233
rect 15292 4224 15344 4276
rect 16028 4224 16080 4276
rect 4068 4156 4120 4208
rect 4160 4088 4212 4140
rect 8392 4156 8444 4208
rect 3516 4020 3568 4072
rect 4068 4020 4120 4072
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 8208 4088 8260 4140
rect 5540 3952 5592 4004
rect 8668 4020 8720 4072
rect 9496 4020 9548 4072
rect 9680 4020 9732 4072
rect 9956 4020 10008 4072
rect 10600 4063 10652 4072
rect 10600 4029 10609 4063
rect 10609 4029 10643 4063
rect 10643 4029 10652 4063
rect 10600 4020 10652 4029
rect 12532 4088 12584 4140
rect 14096 4088 14148 4140
rect 14924 4088 14976 4140
rect 3332 3884 3384 3936
rect 4712 3884 4764 3936
rect 5724 3884 5776 3936
rect 5816 3884 5868 3936
rect 8944 3884 8996 3936
rect 9496 3884 9548 3936
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 15844 4020 15896 4072
rect 16396 4063 16448 4072
rect 16396 4029 16397 4063
rect 16397 4029 16431 4063
rect 16431 4029 16448 4063
rect 16396 4020 16448 4029
rect 13728 3952 13780 4004
rect 14188 3995 14240 4004
rect 14188 3961 14197 3995
rect 14197 3961 14231 3995
rect 14231 3961 14240 3995
rect 14188 3952 14240 3961
rect 12716 3927 12768 3936
rect 12716 3893 12725 3927
rect 12725 3893 12759 3927
rect 12759 3893 12768 3927
rect 12716 3884 12768 3893
rect 15016 3884 15068 3936
rect 15292 3927 15344 3936
rect 15292 3893 15301 3927
rect 15301 3893 15335 3927
rect 15335 3893 15344 3927
rect 15292 3884 15344 3893
rect 16212 3927 16264 3936
rect 16212 3893 16221 3927
rect 16221 3893 16255 3927
rect 16255 3893 16264 3927
rect 16212 3884 16264 3893
rect 6410 3782 6462 3834
rect 6474 3782 6526 3834
rect 6538 3782 6590 3834
rect 6602 3782 6654 3834
rect 11838 3782 11890 3834
rect 11902 3782 11954 3834
rect 11966 3782 12018 3834
rect 12030 3782 12082 3834
rect 2228 3680 2280 3732
rect 4528 3680 4580 3732
rect 5356 3680 5408 3732
rect 3056 3612 3108 3664
rect 8576 3680 8628 3732
rect 9956 3680 10008 3732
rect 6920 3612 6972 3664
rect 8208 3612 8260 3664
rect 9588 3612 9640 3664
rect 10600 3680 10652 3732
rect 12992 3680 13044 3732
rect 13728 3723 13780 3732
rect 13728 3689 13737 3723
rect 13737 3689 13771 3723
rect 13771 3689 13780 3723
rect 13728 3680 13780 3689
rect 3424 3476 3476 3528
rect 8300 3544 8352 3596
rect 5724 3476 5776 3528
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 7748 3476 7800 3528
rect 9956 3544 10008 3596
rect 8576 3476 8628 3528
rect 12532 3612 12584 3664
rect 13360 3612 13412 3664
rect 11428 3587 11480 3596
rect 3056 3340 3108 3392
rect 4252 3408 4304 3460
rect 4528 3408 4580 3460
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 6000 3340 6052 3392
rect 8760 3408 8812 3460
rect 11428 3553 11437 3587
rect 11437 3553 11471 3587
rect 11471 3553 11480 3587
rect 11428 3544 11480 3553
rect 11612 3587 11664 3596
rect 11612 3553 11621 3587
rect 11621 3553 11655 3587
rect 11655 3553 11664 3587
rect 11612 3544 11664 3553
rect 11704 3587 11756 3596
rect 11704 3553 11713 3587
rect 11713 3553 11747 3587
rect 11747 3553 11756 3587
rect 11704 3544 11756 3553
rect 12164 3544 12216 3596
rect 12440 3544 12492 3596
rect 15200 3612 15252 3664
rect 16212 3612 16264 3664
rect 14924 3587 14976 3596
rect 14924 3553 14933 3587
rect 14933 3553 14967 3587
rect 14967 3553 14976 3587
rect 14924 3544 14976 3553
rect 15200 3519 15252 3528
rect 7288 3340 7340 3392
rect 8208 3383 8260 3392
rect 8208 3349 8217 3383
rect 8217 3349 8251 3383
rect 8251 3349 8260 3383
rect 8208 3340 8260 3349
rect 8484 3340 8536 3392
rect 9588 3340 9640 3392
rect 15200 3485 15209 3519
rect 15209 3485 15243 3519
rect 15243 3485 15252 3519
rect 15200 3476 15252 3485
rect 15844 3476 15896 3528
rect 13728 3408 13780 3460
rect 11060 3340 11112 3392
rect 3696 3238 3748 3290
rect 3760 3238 3812 3290
rect 3824 3238 3876 3290
rect 3888 3238 3940 3290
rect 9124 3238 9176 3290
rect 9188 3238 9240 3290
rect 9252 3238 9304 3290
rect 9316 3238 9368 3290
rect 14552 3238 14604 3290
rect 14616 3238 14668 3290
rect 14680 3238 14732 3290
rect 14744 3238 14796 3290
rect 4068 3136 4120 3188
rect 4528 3179 4580 3188
rect 4528 3145 4537 3179
rect 4537 3145 4571 3179
rect 4571 3145 4580 3179
rect 4528 3136 4580 3145
rect 7748 3136 7800 3188
rect 3976 3068 4028 3120
rect 5816 3068 5868 3120
rect 1952 3000 2004 3052
rect 480 2932 532 2984
rect 4528 2932 4580 2984
rect 3332 2864 3384 2916
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 9496 3136 9548 3188
rect 11428 3136 11480 3188
rect 13820 3179 13872 3188
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 14188 3136 14240 3188
rect 15016 3179 15068 3188
rect 15016 3145 15025 3179
rect 15025 3145 15059 3179
rect 15059 3145 15068 3179
rect 15016 3136 15068 3145
rect 15200 3136 15252 3188
rect 11244 3000 11296 3052
rect 5448 2864 5500 2916
rect 8208 2864 8260 2916
rect 9680 2864 9732 2916
rect 10600 2864 10652 2916
rect 4620 2796 4672 2848
rect 4712 2839 4764 2848
rect 4712 2805 4721 2839
rect 4721 2805 4755 2839
rect 4755 2805 4764 2839
rect 4712 2796 4764 2805
rect 5172 2796 5224 2848
rect 15568 3068 15620 3120
rect 11704 3000 11756 3052
rect 15016 3000 15068 3052
rect 12256 2975 12308 2984
rect 12256 2941 12262 2975
rect 12262 2941 12296 2975
rect 12296 2941 12308 2975
rect 12256 2932 12308 2941
rect 12164 2796 12216 2848
rect 13360 2975 13412 2984
rect 13360 2941 13369 2975
rect 13369 2941 13403 2975
rect 13403 2941 13412 2975
rect 13360 2932 13412 2941
rect 14280 2932 14332 2984
rect 15844 2975 15896 2984
rect 15844 2941 15853 2975
rect 15853 2941 15887 2975
rect 15887 2941 15896 2975
rect 15844 2932 15896 2941
rect 16028 2932 16080 2984
rect 15476 2864 15528 2916
rect 13176 2839 13228 2848
rect 13176 2805 13185 2839
rect 13185 2805 13219 2839
rect 13219 2805 13228 2839
rect 13176 2796 13228 2805
rect 15016 2796 15068 2848
rect 6410 2694 6462 2746
rect 6474 2694 6526 2746
rect 6538 2694 6590 2746
rect 6602 2694 6654 2746
rect 11838 2694 11890 2746
rect 11902 2694 11954 2746
rect 11966 2694 12018 2746
rect 12030 2694 12082 2746
rect 3424 2592 3476 2644
rect 1860 2456 1912 2508
rect 4160 2524 4212 2576
rect 4620 2592 4672 2644
rect 5632 2592 5684 2644
rect 6000 2592 6052 2644
rect 4528 2567 4580 2576
rect 4252 2499 4304 2508
rect 4252 2465 4261 2499
rect 4261 2465 4295 2499
rect 4295 2465 4304 2499
rect 4252 2456 4304 2465
rect 4528 2533 4537 2567
rect 4537 2533 4571 2567
rect 4571 2533 4580 2567
rect 4528 2524 4580 2533
rect 5724 2524 5776 2576
rect 7380 2592 7432 2644
rect 9680 2592 9732 2644
rect 10600 2592 10652 2644
rect 11428 2592 11480 2644
rect 12256 2635 12308 2644
rect 12256 2601 12265 2635
rect 12265 2601 12299 2635
rect 12299 2601 12308 2635
rect 12256 2592 12308 2601
rect 15476 2635 15528 2644
rect 15476 2601 15485 2635
rect 15485 2601 15519 2635
rect 15519 2601 15528 2635
rect 15476 2592 15528 2601
rect 4712 2456 4764 2508
rect 6000 2499 6052 2508
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 4804 2388 4856 2440
rect 4344 2320 4396 2372
rect 5448 2388 5500 2440
rect 5356 2363 5408 2372
rect 5356 2329 5365 2363
rect 5365 2329 5399 2363
rect 5399 2329 5408 2363
rect 8576 2456 8628 2508
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 11060 2524 11112 2576
rect 13176 2524 13228 2576
rect 13728 2567 13780 2576
rect 13728 2533 13737 2567
rect 13737 2533 13771 2567
rect 13771 2533 13780 2567
rect 13728 2524 13780 2533
rect 15568 2524 15620 2576
rect 11612 2456 11664 2508
rect 14096 2456 14148 2508
rect 15660 2499 15712 2508
rect 15660 2465 15669 2499
rect 15669 2465 15703 2499
rect 15703 2465 15712 2499
rect 15660 2456 15712 2465
rect 17500 2456 17552 2508
rect 5356 2320 5408 2329
rect 5632 2252 5684 2304
rect 11428 2320 11480 2372
rect 12716 2320 12768 2372
rect 16488 2295 16540 2304
rect 16488 2261 16497 2295
rect 16497 2261 16531 2295
rect 16531 2261 16540 2295
rect 16488 2252 16540 2261
rect 3696 2150 3748 2202
rect 3760 2150 3812 2202
rect 3824 2150 3876 2202
rect 3888 2150 3940 2202
rect 9124 2150 9176 2202
rect 9188 2150 9240 2202
rect 9252 2150 9304 2202
rect 9316 2150 9368 2202
rect 14552 2150 14604 2202
rect 14616 2150 14668 2202
rect 14680 2150 14732 2202
rect 14744 2150 14796 2202
rect 4436 2048 4488 2100
rect 16488 2048 16540 2100
<< metal2 >>
rect 938 19892 994 20692
rect 2318 19892 2374 20692
rect 4158 19892 4214 20692
rect 5998 19892 6054 20692
rect 7838 19892 7894 20692
rect 9678 19892 9734 20692
rect 11058 19892 11114 20692
rect 12898 19892 12954 20692
rect 14738 19892 14794 20692
rect 16578 19892 16634 20692
rect 17958 19892 18014 20692
rect 952 18290 980 19892
rect 1766 18456 1822 18465
rect 1766 18391 1822 18400
rect 940 18284 992 18290
rect 940 18226 992 18232
rect 1780 18222 1808 18391
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 2332 18170 2360 19892
rect 3670 18524 3966 18544
rect 3726 18522 3750 18524
rect 3806 18522 3830 18524
rect 3886 18522 3910 18524
rect 3748 18470 3750 18522
rect 3812 18470 3824 18522
rect 3886 18470 3888 18522
rect 3726 18468 3750 18470
rect 3806 18468 3830 18470
rect 3886 18468 3910 18470
rect 3670 18448 3966 18468
rect 4172 18306 4200 19892
rect 4080 18278 4200 18306
rect 4080 18222 4108 18278
rect 4068 18216 4120 18222
rect 2332 18142 2452 18170
rect 4068 18158 4120 18164
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 1964 17814 1992 18022
rect 1952 17808 2004 17814
rect 1952 17750 2004 17756
rect 2332 17746 2360 18022
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2424 17134 2452 18142
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 1492 16516 1544 16522
rect 1492 16458 1544 16464
rect 1504 16114 1532 16458
rect 2516 16114 2544 17478
rect 3344 17338 3372 17478
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2608 16250 2636 16390
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 1400 13456 1452 13462
rect 1400 13398 1452 13404
rect 1412 12442 1440 13398
rect 1504 12850 1532 16050
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1688 15162 1716 15982
rect 2608 15910 2636 16186
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 1950 15736 2006 15745
rect 1950 15671 2006 15680
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1872 14618 1900 15302
rect 1964 14958 1992 15671
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 2056 14482 2084 15846
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2240 14822 2268 15438
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2240 14550 2268 14758
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2688 13728 2740 13734
rect 2688 13670 2740 13676
rect 2700 13462 2728 13670
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2778 13016 2834 13025
rect 2778 12951 2834 12960
rect 1492 12844 1544 12850
rect 1492 12786 1544 12792
rect 2792 12782 2820 12951
rect 2884 12850 2912 16934
rect 3252 16590 3280 16934
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3252 15978 3280 16526
rect 3344 16454 3372 16730
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3344 16046 3372 16390
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3240 15972 3292 15978
rect 3240 15914 3292 15920
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2976 14482 3004 15506
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2976 13530 3004 14418
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 1400 12436 1452 12442
rect 1400 12378 1452 12384
rect 1872 12306 1900 12582
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2148 11354 2176 12242
rect 2976 12238 3004 13126
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 3068 12374 3096 12650
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1780 10985 1808 11154
rect 1766 10976 1822 10985
rect 1766 10911 1822 10920
rect 2148 10606 2176 11290
rect 2240 10606 2268 12174
rect 2976 11762 3004 12174
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2332 10538 2360 11154
rect 2424 11014 2452 11290
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2424 10606 2452 10950
rect 2608 10810 2636 11562
rect 2688 11552 2740 11558
rect 2688 11494 2740 11500
rect 2700 11218 2728 11494
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2320 10532 2372 10538
rect 2320 10474 2372 10480
rect 1400 10192 1452 10198
rect 1400 10134 1452 10140
rect 1412 9178 1440 10134
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1872 8922 1900 8978
rect 2044 8968 2096 8974
rect 1872 8916 2044 8922
rect 1872 8910 2096 8916
rect 1872 8894 2084 8910
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 8090 1716 8366
rect 2056 8294 2084 8894
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2044 8288 2096 8294
rect 1950 8256 2006 8265
rect 2044 8230 2096 8236
rect 1950 8191 2006 8200
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1964 7954 1992 8191
rect 2332 7954 2360 8774
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2424 7834 2452 10542
rect 2976 10062 3004 11698
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 3068 10198 3096 10406
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 3252 9518 3280 10542
rect 3344 10266 3372 15982
rect 3528 14006 3556 17614
rect 3670 17436 3966 17456
rect 3726 17434 3750 17436
rect 3806 17434 3830 17436
rect 3886 17434 3910 17436
rect 3748 17382 3750 17434
rect 3812 17382 3824 17434
rect 3886 17382 3888 17434
rect 3726 17380 3750 17382
rect 3806 17380 3830 17382
rect 3886 17380 3910 17382
rect 3670 17360 3966 17380
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 4528 17060 4580 17066
rect 4528 17002 4580 17008
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 3670 16348 3966 16368
rect 3726 16346 3750 16348
rect 3806 16346 3830 16348
rect 3886 16346 3910 16348
rect 3748 16294 3750 16346
rect 3812 16294 3824 16346
rect 3886 16294 3888 16346
rect 3726 16292 3750 16294
rect 3806 16292 3830 16294
rect 3886 16292 3910 16294
rect 3670 16272 3966 16292
rect 3670 15260 3966 15280
rect 3726 15258 3750 15260
rect 3806 15258 3830 15260
rect 3886 15258 3910 15260
rect 3748 15206 3750 15258
rect 3812 15206 3824 15258
rect 3886 15206 3888 15258
rect 3726 15204 3750 15206
rect 3806 15204 3830 15206
rect 3886 15204 3910 15206
rect 3670 15184 3966 15204
rect 4172 15162 4200 16594
rect 4448 16250 4476 17002
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4436 15972 4488 15978
rect 4436 15914 4488 15920
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 3976 14952 4028 14958
rect 4172 14940 4200 15098
rect 4028 14912 4200 14940
rect 4344 14952 4396 14958
rect 3976 14894 4028 14900
rect 4344 14894 4396 14900
rect 3700 14884 3752 14890
rect 3700 14826 3752 14832
rect 3712 14618 3740 14826
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3988 14482 4016 14894
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3670 14172 3966 14192
rect 3726 14170 3750 14172
rect 3806 14170 3830 14172
rect 3886 14170 3910 14172
rect 3748 14118 3750 14170
rect 3812 14118 3824 14170
rect 3886 14118 3888 14170
rect 3726 14116 3750 14118
rect 3806 14116 3830 14118
rect 3886 14116 3910 14118
rect 3670 14096 3966 14116
rect 4356 14006 4384 14894
rect 4448 14550 4476 15914
rect 4540 15910 4568 17002
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4632 15570 4660 15982
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4632 14550 4660 15302
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 4172 13818 4200 13874
rect 4356 13818 4384 13942
rect 3528 12306 3556 13806
rect 4172 13790 4384 13818
rect 4436 13864 4488 13870
rect 4436 13806 4488 13812
rect 3670 13084 3966 13104
rect 3726 13082 3750 13084
rect 3806 13082 3830 13084
rect 3886 13082 3910 13084
rect 3748 13030 3750 13082
rect 3812 13030 3824 13082
rect 3886 13030 3888 13082
rect 3726 13028 3750 13030
rect 3806 13028 3830 13030
rect 3886 13028 3910 13030
rect 3670 13008 3966 13028
rect 4172 12782 4200 13790
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3528 12102 3556 12242
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3670 11996 3966 12016
rect 3726 11994 3750 11996
rect 3806 11994 3830 11996
rect 3886 11994 3910 11996
rect 3748 11942 3750 11994
rect 3812 11942 3824 11994
rect 3886 11942 3888 11994
rect 3726 11940 3750 11942
rect 3806 11940 3830 11942
rect 3886 11940 3910 11942
rect 3670 11920 3966 11940
rect 4080 11694 4108 12582
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3670 10908 3966 10928
rect 3726 10906 3750 10908
rect 3806 10906 3830 10908
rect 3886 10906 3910 10908
rect 3748 10854 3750 10906
rect 3812 10854 3824 10906
rect 3886 10854 3888 10906
rect 3726 10852 3750 10854
rect 3806 10852 3830 10854
rect 3886 10852 3910 10854
rect 3670 10832 3966 10852
rect 4080 10810 4108 11086
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3670 9820 3966 9840
rect 3726 9818 3750 9820
rect 3806 9818 3830 9820
rect 3886 9818 3910 9820
rect 3748 9766 3750 9818
rect 3812 9766 3824 9818
rect 3886 9766 3888 9818
rect 3726 9764 3750 9766
rect 3806 9764 3830 9766
rect 3886 9764 3910 9766
rect 3670 9744 3966 9764
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2608 8634 2636 8978
rect 2700 8838 2728 9114
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2516 7954 2544 8230
rect 2608 8022 2636 8570
rect 2596 8016 2648 8022
rect 2596 7958 2648 7964
rect 2700 7954 2728 8774
rect 3528 8362 3556 9318
rect 3670 8732 3966 8752
rect 3726 8730 3750 8732
rect 3806 8730 3830 8732
rect 3886 8730 3910 8732
rect 3748 8678 3750 8730
rect 3812 8678 3824 8730
rect 3886 8678 3888 8730
rect 3726 8676 3750 8678
rect 3806 8676 3830 8678
rect 3886 8676 3910 8678
rect 3670 8656 3966 8676
rect 4356 8362 4384 12038
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4080 8090 4108 8298
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2332 7806 2452 7834
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 6934 1716 7142
rect 1676 6928 1728 6934
rect 1676 6870 1728 6876
rect 2332 6798 2360 7806
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 3670 7644 3966 7664
rect 3726 7642 3750 7644
rect 3806 7642 3830 7644
rect 3886 7642 3910 7644
rect 3748 7590 3750 7642
rect 3812 7590 3824 7642
rect 3886 7590 3888 7642
rect 3726 7588 3750 7590
rect 3806 7588 3830 7590
rect 3886 7588 3910 7590
rect 3670 7568 3966 7588
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2044 6792 2096 6798
rect 1964 6752 2044 6780
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5914 1624 6054
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5545 1440 5714
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1964 5166 1992 6752
rect 2044 6734 2096 6740
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2424 6458 2452 6870
rect 3160 6458 3188 7278
rect 3528 7206 3556 7482
rect 4080 7342 4108 7482
rect 4264 7410 4292 7686
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 1964 4622 1992 5102
rect 2228 5092 2280 5098
rect 2228 5034 2280 5040
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1964 3058 1992 4558
rect 2240 3738 2268 5034
rect 2792 4690 2820 6190
rect 3528 5370 3556 7142
rect 3670 6556 3966 6576
rect 3726 6554 3750 6556
rect 3806 6554 3830 6556
rect 3886 6554 3910 6556
rect 3748 6502 3750 6554
rect 3812 6502 3824 6554
rect 3886 6502 3888 6554
rect 3726 6500 3750 6502
rect 3806 6500 3830 6502
rect 3886 6500 3910 6502
rect 3670 6480 3966 6500
rect 4264 6322 4292 7142
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4172 5914 4200 6122
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 3670 5468 3966 5488
rect 3726 5466 3750 5468
rect 3806 5466 3830 5468
rect 3886 5466 3910 5468
rect 3748 5414 3750 5466
rect 3812 5414 3824 5466
rect 3886 5414 3888 5466
rect 3726 5412 3750 5414
rect 3806 5412 3830 5414
rect 3886 5412 3910 5414
rect 3670 5392 3966 5412
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2976 4826 3004 5034
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 4080 4690 4108 5714
rect 4356 5166 4384 8298
rect 4344 5160 4396 5166
rect 4344 5102 4396 5108
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4080 4486 4108 4626
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3670 4380 3966 4400
rect 3726 4378 3750 4380
rect 3806 4378 3830 4380
rect 3886 4378 3910 4380
rect 3748 4326 3750 4378
rect 3812 4326 3824 4378
rect 3886 4326 3888 4378
rect 3726 4324 3750 4326
rect 3806 4324 3830 4326
rect 3886 4324 3910 4326
rect 3670 4304 3966 4324
rect 4080 4214 4108 4422
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 3068 3398 3096 3606
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 492 800 520 2926
rect 3344 2922 3372 3878
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3332 2916 3384 2922
rect 3332 2858 3384 2864
rect 3436 2650 3464 3470
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 1872 800 1900 2450
rect 3528 1442 3556 4014
rect 3670 3292 3966 3312
rect 3726 3290 3750 3292
rect 3806 3290 3830 3292
rect 3886 3290 3910 3292
rect 3748 3238 3750 3290
rect 3812 3238 3824 3290
rect 3886 3238 3888 3290
rect 3726 3236 3750 3238
rect 3806 3236 3830 3238
rect 3886 3236 3910 3238
rect 3670 3216 3966 3236
rect 4080 3194 4108 4014
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 3988 2825 4016 3062
rect 3974 2816 4030 2825
rect 3974 2751 4030 2760
rect 4172 2582 4200 4082
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4264 2514 4292 3402
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 4356 2378 4384 5102
rect 4344 2372 4396 2378
rect 4344 2314 4396 2320
rect 3670 2204 3966 2224
rect 3726 2202 3750 2204
rect 3806 2202 3830 2204
rect 3886 2202 3910 2204
rect 3748 2150 3750 2202
rect 3812 2150 3824 2202
rect 3886 2150 3888 2202
rect 3726 2148 3750 2150
rect 3806 2148 3830 2150
rect 3886 2148 3910 2150
rect 3670 2128 3966 2148
rect 4448 2106 4476 13806
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4528 12912 4580 12918
rect 4528 12854 4580 12860
rect 4540 11762 4568 12854
rect 4632 11898 4660 12922
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4632 11558 4660 11834
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4724 10146 4752 18022
rect 4816 17542 4844 18158
rect 5092 17678 5120 18158
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 5092 17202 5120 17614
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 5276 17134 5304 18090
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 5368 17134 5396 17478
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 4816 16658 4844 17070
rect 5552 17066 5580 18158
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 16726 5212 16934
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 5552 15706 5580 17002
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 5920 16250 5948 16662
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 6012 15570 6040 19892
rect 7852 18358 7880 19892
rect 9098 18524 9394 18544
rect 9154 18522 9178 18524
rect 9234 18522 9258 18524
rect 9314 18522 9338 18524
rect 9176 18470 9178 18522
rect 9240 18470 9252 18522
rect 9314 18470 9316 18522
rect 9154 18468 9178 18470
rect 9234 18468 9258 18470
rect 9314 18468 9338 18470
rect 9098 18448 9394 18468
rect 7840 18352 7892 18358
rect 7840 18294 7892 18300
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6104 17814 6132 18022
rect 6384 17980 6680 18000
rect 6440 17978 6464 17980
rect 6520 17978 6544 17980
rect 6600 17978 6624 17980
rect 6462 17926 6464 17978
rect 6526 17926 6538 17978
rect 6600 17926 6602 17978
rect 6440 17924 6464 17926
rect 6520 17924 6544 17926
rect 6600 17924 6624 17926
rect 6384 17904 6680 17924
rect 6840 17882 6868 18022
rect 8588 17882 8616 18090
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 6092 17808 6144 17814
rect 6092 17750 6144 17756
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 6748 17270 6776 17614
rect 7116 17338 7144 17614
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 6736 17264 6788 17270
rect 6736 17206 6788 17212
rect 6384 16892 6680 16912
rect 6440 16890 6464 16892
rect 6520 16890 6544 16892
rect 6600 16890 6624 16892
rect 6462 16838 6464 16890
rect 6526 16838 6538 16890
rect 6600 16838 6602 16890
rect 6440 16836 6464 16838
rect 6520 16836 6544 16838
rect 6600 16836 6624 16838
rect 6384 16816 6680 16836
rect 6384 15804 6680 15824
rect 6440 15802 6464 15804
rect 6520 15802 6544 15804
rect 6600 15802 6624 15804
rect 6462 15750 6464 15802
rect 6526 15750 6538 15802
rect 6600 15750 6602 15802
rect 6440 15748 6464 15750
rect 6520 15748 6544 15750
rect 6600 15748 6624 15750
rect 6384 15728 6680 15748
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 6748 15366 6776 17206
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7668 16998 7696 17138
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7116 15570 7144 15846
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6748 15162 6776 15302
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5552 14414 5580 15030
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 14074 5580 14350
rect 5736 14074 5764 14826
rect 5828 14822 5856 14894
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 5828 14618 5856 14758
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 6012 14278 6040 14758
rect 6384 14716 6680 14736
rect 6440 14714 6464 14716
rect 6520 14714 6544 14716
rect 6600 14714 6624 14716
rect 6462 14662 6464 14714
rect 6526 14662 6538 14714
rect 6600 14662 6602 14714
rect 6440 14660 6464 14662
rect 6520 14660 6544 14662
rect 6600 14660 6624 14662
rect 6384 14640 6680 14660
rect 6748 14550 6776 14894
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5552 13734 5580 14010
rect 6656 13870 6684 14418
rect 6748 14074 6776 14486
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 6384 13628 6680 13648
rect 6440 13626 6464 13628
rect 6520 13626 6544 13628
rect 6600 13626 6624 13628
rect 6462 13574 6464 13626
rect 6526 13574 6538 13626
rect 6600 13574 6602 13626
rect 6440 13572 6464 13574
rect 6520 13572 6544 13574
rect 6600 13572 6624 13574
rect 6384 13552 6680 13572
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4816 12374 4844 13126
rect 5000 12918 5028 13330
rect 5184 12986 5212 13330
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 5276 12782 5304 13262
rect 5552 12782 5580 13398
rect 6840 13190 6868 15506
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7024 13938 7052 14214
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7116 13394 7144 15506
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5276 12646 5304 12718
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 11286 5120 11494
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 5276 10810 5304 12582
rect 5552 12442 5580 12718
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5828 12238 5856 12582
rect 5920 12306 5948 13126
rect 6012 12782 6040 13126
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 6384 12540 6680 12560
rect 6440 12538 6464 12540
rect 6520 12538 6544 12540
rect 6600 12538 6624 12540
rect 6462 12486 6464 12538
rect 6526 12486 6538 12538
rect 6600 12486 6602 12538
rect 6440 12484 6464 12486
rect 6520 12484 6544 12486
rect 6600 12484 6624 12486
rect 6384 12464 6680 12484
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5552 11150 5580 12174
rect 6384 11452 6680 11472
rect 6440 11450 6464 11452
rect 6520 11450 6544 11452
rect 6600 11450 6624 11452
rect 6462 11398 6464 11450
rect 6526 11398 6538 11450
rect 6600 11398 6602 11450
rect 6440 11396 6464 11398
rect 6520 11396 6544 11398
rect 6600 11396 6624 11398
rect 6384 11376 6680 11396
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5092 10266 5120 10542
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4632 10118 4752 10146
rect 4632 8022 4660 10118
rect 4710 9616 4766 9625
rect 4710 9551 4766 9560
rect 4724 9518 4752 9551
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 5264 9512 5316 9518
rect 5316 9472 5396 9500
rect 5264 9454 5316 9460
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 9110 4752 9318
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4724 8362 4752 8502
rect 5368 8362 5396 9472
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5460 8430 5488 8502
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5368 8090 5396 8298
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4540 5370 4568 7890
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4540 3738 4568 4558
rect 4724 3942 4752 7890
rect 5460 7886 5488 8366
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5460 7546 5488 7822
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 4816 6934 4844 7142
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 6254 4936 6734
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 4908 5914 4936 6190
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4816 4570 4844 5306
rect 4908 4826 4936 5850
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4896 4616 4948 4622
rect 4816 4564 4896 4570
rect 4816 4558 4948 4564
rect 4816 4542 4936 4558
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4528 3460 4580 3466
rect 4528 3402 4580 3408
rect 4540 3194 4568 3402
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4540 2582 4568 2926
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4632 2650 4660 2790
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 4724 2514 4752 2790
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 4816 2446 4844 4542
rect 5184 4078 5212 6190
rect 5460 5370 5488 7142
rect 5644 6254 5672 11290
rect 5816 11280 5868 11286
rect 5816 11222 5868 11228
rect 5828 10266 5856 11222
rect 6384 10364 6680 10384
rect 6440 10362 6464 10364
rect 6520 10362 6544 10364
rect 6600 10362 6624 10364
rect 6462 10310 6464 10362
rect 6526 10310 6538 10362
rect 6600 10310 6602 10362
rect 6440 10308 6464 10310
rect 6520 10308 6544 10310
rect 6600 10308 6624 10310
rect 6384 10288 6680 10308
rect 6932 10266 6960 12310
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7024 10266 7052 10950
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7116 10198 7144 10950
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7208 9654 7236 16730
rect 7668 16658 7696 16934
rect 7852 16658 7880 17070
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 7944 16726 7972 16934
rect 8220 16794 8248 17002
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7668 16250 7696 16594
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7944 16114 7972 16662
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 8220 16046 8248 16594
rect 8772 16250 8800 17750
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8956 16046 8984 18158
rect 9098 17436 9394 17456
rect 9154 17434 9178 17436
rect 9234 17434 9258 17436
rect 9314 17434 9338 17436
rect 9176 17382 9178 17434
rect 9240 17382 9252 17434
rect 9314 17382 9316 17434
rect 9154 17380 9178 17382
rect 9234 17380 9258 17382
rect 9314 17380 9338 17382
rect 9098 17360 9394 17380
rect 9496 17060 9548 17066
rect 9496 17002 9548 17008
rect 9098 16348 9394 16368
rect 9154 16346 9178 16348
rect 9234 16346 9258 16348
rect 9314 16346 9338 16348
rect 9176 16294 9178 16346
rect 9240 16294 9252 16346
rect 9314 16294 9316 16346
rect 9154 16292 9178 16294
rect 9234 16292 9258 16294
rect 9314 16292 9338 16294
rect 9098 16272 9394 16292
rect 9508 16250 9536 17002
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 8220 15910 8248 15982
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7576 14890 7604 15302
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 8128 14550 8156 15506
rect 8220 15162 8248 15846
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8956 14618 8984 15982
rect 9692 15978 9720 19892
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9784 16794 9812 17614
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9876 16182 9904 18158
rect 10048 17808 10100 17814
rect 10048 17750 10100 17756
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9876 15570 9904 15846
rect 9968 15638 9996 16594
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9098 15260 9394 15280
rect 9154 15258 9178 15260
rect 9234 15258 9258 15260
rect 9314 15258 9338 15260
rect 9176 15206 9178 15258
rect 9240 15206 9252 15258
rect 9314 15206 9316 15258
rect 9154 15204 9178 15206
rect 9234 15204 9258 15206
rect 9314 15204 9338 15206
rect 9098 15184 9394 15204
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8116 14544 8168 14550
rect 8956 14498 8984 14554
rect 8116 14486 8168 14492
rect 8864 14470 8984 14498
rect 9496 14476 9548 14482
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7300 13530 7328 13738
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 6288 8974 6316 9590
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6384 9276 6680 9296
rect 6440 9274 6464 9276
rect 6520 9274 6544 9276
rect 6600 9274 6624 9276
rect 6462 9222 6464 9274
rect 6526 9222 6538 9274
rect 6600 9222 6602 9274
rect 6440 9220 6464 9222
rect 6520 9220 6544 9222
rect 6600 9220 6624 9222
rect 6384 9200 6680 9220
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6288 8634 6316 8910
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5828 7478 5856 8366
rect 6288 8294 6316 8570
rect 6840 8430 6868 9318
rect 7116 9178 7144 9454
rect 7208 9382 7236 9590
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7116 8430 7144 9114
rect 7208 8430 7236 9318
rect 7300 8498 7328 12650
rect 7576 11694 7604 13262
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7852 12986 7880 13194
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7944 12714 7972 13262
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8588 12782 8616 13126
rect 8680 12986 8708 13126
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8680 12714 8708 12922
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7760 11898 7788 12310
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 10470 7420 11086
rect 7484 11082 7512 11290
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7392 10198 7420 10406
rect 7484 10266 7512 11018
rect 7576 11014 7604 11630
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 9178 7512 9454
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7392 8634 7420 8910
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6384 8188 6680 8208
rect 6440 8186 6464 8188
rect 6520 8186 6544 8188
rect 6600 8186 6624 8188
rect 6462 8134 6464 8186
rect 6526 8134 6538 8186
rect 6600 8134 6602 8186
rect 6440 8132 6464 8134
rect 6520 8132 6544 8134
rect 6600 8132 6624 8134
rect 6384 8112 6680 8132
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5736 6118 5764 7346
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5736 5302 5764 6054
rect 5828 5778 5856 7414
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 6934 6132 7142
rect 6384 7100 6680 7120
rect 6440 7098 6464 7100
rect 6520 7098 6544 7100
rect 6600 7098 6624 7100
rect 6462 7046 6464 7098
rect 6526 7046 6538 7098
rect 6600 7046 6602 7098
rect 6440 7044 6464 7046
rect 6520 7044 6544 7046
rect 6600 7044 6624 7046
rect 6384 7024 6680 7044
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6748 6866 6776 8230
rect 7852 8022 7880 8978
rect 8036 8838 8064 12582
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8404 10538 8432 11018
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8128 8634 8156 10066
rect 8496 9994 8524 12650
rect 8772 12594 8800 13806
rect 8864 12730 8892 14470
rect 9496 14418 9548 14424
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8956 13870 8984 14282
rect 9098 14172 9394 14192
rect 9154 14170 9178 14172
rect 9234 14170 9258 14172
rect 9314 14170 9338 14172
rect 9176 14118 9178 14170
rect 9240 14118 9252 14170
rect 9314 14118 9316 14170
rect 9154 14116 9178 14118
rect 9234 14116 9258 14118
rect 9314 14116 9338 14118
rect 9098 14096 9394 14116
rect 9508 14074 9536 14418
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9692 14006 9720 14962
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9784 14618 9812 14826
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 10060 14074 10088 17750
rect 10152 17202 10180 18226
rect 11072 18154 11100 19892
rect 12912 18290 12940 19892
rect 14752 18714 14780 19892
rect 14384 18686 14780 18714
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 11812 17980 12108 18000
rect 11868 17978 11892 17980
rect 11948 17978 11972 17980
rect 12028 17978 12052 17980
rect 11890 17926 11892 17978
rect 11954 17926 11966 17978
rect 12028 17926 12030 17978
rect 11868 17924 11892 17926
rect 11948 17924 11972 17926
rect 12028 17924 12052 17926
rect 11812 17904 12108 17924
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 10152 16454 10180 17138
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10428 16454 10456 16730
rect 10520 16658 10548 16934
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 15910 10456 16390
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10612 15570 10640 15846
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10612 15162 10640 15506
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10704 14550 10732 16594
rect 10888 15570 10916 17478
rect 11812 16892 12108 16912
rect 11868 16890 11892 16892
rect 11948 16890 11972 16892
rect 12028 16890 12052 16892
rect 11890 16838 11892 16890
rect 11954 16838 11966 16890
rect 12028 16838 12030 16890
rect 11868 16836 11892 16838
rect 11948 16836 11972 16838
rect 12028 16836 12052 16838
rect 11812 16816 12108 16836
rect 12072 16516 12124 16522
rect 12072 16458 12124 16464
rect 12084 16046 12112 16458
rect 12176 16046 12204 18226
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12360 18086 12388 18158
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12268 16658 12296 16934
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 12268 15994 12296 16594
rect 12360 16522 12388 18022
rect 12912 17678 12940 18022
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12452 16794 12480 17478
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 13188 16794 13216 17002
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 12452 16590 12480 16730
rect 13372 16726 13400 18022
rect 13636 17808 13688 17814
rect 13636 17750 13688 17756
rect 13818 17776 13874 17785
rect 13648 16794 13676 17750
rect 13818 17711 13874 17720
rect 13728 17060 13780 17066
rect 13728 17002 13780 17008
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12452 16046 12480 16526
rect 13280 16046 13308 16594
rect 13740 16250 13768 17002
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 12440 16040 12492 16046
rect 11256 15706 11284 15982
rect 12268 15978 12388 15994
rect 12440 15982 12492 15988
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 12268 15972 12400 15978
rect 12268 15966 12348 15972
rect 12348 15914 12400 15920
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 11812 15804 12108 15824
rect 11868 15802 11892 15804
rect 11948 15802 11972 15804
rect 12028 15802 12052 15804
rect 11890 15750 11892 15802
rect 11954 15750 11966 15802
rect 12028 15750 12030 15802
rect 11868 15748 11892 15750
rect 11948 15748 11972 15750
rect 12028 15748 12052 15750
rect 11812 15728 12108 15748
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10888 15162 10916 15506
rect 11256 15502 11284 15642
rect 12728 15638 12756 15846
rect 13280 15706 13308 15982
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10888 15026 10916 15098
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10692 14544 10744 14550
rect 10692 14486 10744 14492
rect 10888 14482 10916 14962
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10600 14340 10652 14346
rect 10600 14282 10652 14288
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9098 13084 9394 13104
rect 9154 13082 9178 13084
rect 9234 13082 9258 13084
rect 9314 13082 9338 13084
rect 9176 13030 9178 13082
rect 9240 13030 9252 13082
rect 9314 13030 9316 13082
rect 9154 13028 9178 13030
rect 9234 13028 9258 13030
rect 9314 13028 9338 13030
rect 9098 13008 9394 13028
rect 9404 12776 9456 12782
rect 8864 12702 8984 12730
rect 9404 12718 9456 12724
rect 8680 12566 8800 12594
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8588 9625 8616 11154
rect 8574 9616 8630 9625
rect 8574 9551 8630 9560
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7656 7472 7708 7478
rect 7656 7414 7708 7420
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7024 7002 7052 7278
rect 7668 7206 7696 7414
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 7024 6882 7052 6938
rect 6736 6860 6788 6866
rect 7024 6854 7144 6882
rect 6736 6802 6788 6808
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7024 6458 7052 6734
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7116 6254 7144 6854
rect 7668 6662 7696 7142
rect 8220 6798 8248 7278
rect 8496 7206 8524 7414
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7668 6254 7696 6598
rect 8220 6254 8248 6734
rect 8496 6254 8524 7142
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6384 6012 6680 6032
rect 6440 6010 6464 6012
rect 6520 6010 6544 6012
rect 6600 6010 6624 6012
rect 6462 5958 6464 6010
rect 6526 5958 6538 6010
rect 6600 5958 6602 6010
rect 6440 5956 6464 5958
rect 6520 5956 6544 5958
rect 6600 5956 6624 5958
rect 6384 5936 6680 5956
rect 6932 5846 6960 6054
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5920 5166 5948 5510
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 6012 5030 6040 5170
rect 6104 5030 6132 5306
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6012 4826 6040 4966
rect 6384 4924 6680 4944
rect 6440 4922 6464 4924
rect 6520 4922 6544 4924
rect 6600 4922 6624 4924
rect 6462 4870 6464 4922
rect 6526 4870 6538 4922
rect 6600 4870 6602 4922
rect 6440 4868 6464 4870
rect 6520 4868 6544 4870
rect 6600 4868 6624 4870
rect 6384 4848 6680 4868
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 7116 4690 7144 6190
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7392 5370 7420 5646
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7760 5166 7788 5646
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 5644 4282 5672 4626
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5184 2854 5212 4014
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5368 3398 5396 3674
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 5368 2378 5396 3334
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 5460 2446 5488 2858
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5356 2372 5408 2378
rect 5356 2314 5408 2320
rect 4436 2100 4488 2106
rect 4436 2042 4488 2048
rect 3528 1414 3740 1442
rect 3712 800 3740 1414
rect 5552 800 5580 3946
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5736 3534 5764 3878
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5644 2310 5672 2586
rect 5736 2582 5764 3470
rect 5828 3126 5856 3878
rect 6384 3836 6680 3856
rect 6440 3834 6464 3836
rect 6520 3834 6544 3836
rect 6600 3834 6624 3836
rect 6462 3782 6464 3834
rect 6526 3782 6538 3834
rect 6600 3782 6602 3834
rect 6440 3780 6464 3782
rect 6520 3780 6544 3782
rect 6600 3780 6624 3782
rect 6384 3760 6680 3780
rect 6932 3670 6960 4422
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 7760 3534 7788 5102
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 8036 4282 8064 4490
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8220 4146 8248 5510
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8220 3670 8248 4082
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8312 3602 8340 4558
rect 8404 4214 8432 4626
rect 8496 4282 8524 5034
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8392 4208 8444 4214
rect 8392 4150 8444 4156
rect 8588 3738 8616 8298
rect 8680 5846 8708 12566
rect 8956 12458 8984 12702
rect 8772 12430 8984 12458
rect 8772 8498 8800 12430
rect 9416 12186 9444 12718
rect 9508 12306 9536 13126
rect 9600 12442 9628 13874
rect 10612 13802 10640 14282
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10060 13190 10088 13466
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9416 12158 9536 12186
rect 9098 11996 9394 12016
rect 9154 11994 9178 11996
rect 9234 11994 9258 11996
rect 9314 11994 9338 11996
rect 9176 11942 9178 11994
rect 9240 11942 9252 11994
rect 9314 11942 9316 11994
rect 9154 11940 9178 11942
rect 9234 11940 9258 11942
rect 9314 11940 9338 11942
rect 9098 11920 9394 11940
rect 9508 11762 9536 12158
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9098 10908 9394 10928
rect 9154 10906 9178 10908
rect 9234 10906 9258 10908
rect 9314 10906 9338 10908
rect 9176 10854 9178 10906
rect 9240 10854 9252 10906
rect 9314 10854 9316 10906
rect 9154 10852 9178 10854
rect 9234 10852 9258 10854
rect 9314 10852 9338 10854
rect 9098 10832 9394 10852
rect 9508 10606 9536 11698
rect 9600 11286 9628 12378
rect 9692 12170 9720 12650
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9784 11914 9812 12786
rect 10060 12434 10088 13126
rect 10152 12986 10180 13262
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 9876 12406 10088 12434
rect 9876 12306 9904 12406
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9876 12102 9904 12242
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9968 11914 9996 12310
rect 10152 12238 10180 12922
rect 10428 12714 10456 13670
rect 10612 13394 10640 13738
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10612 12374 10640 13330
rect 11164 13258 11192 13806
rect 11348 13734 11376 14894
rect 11812 14716 12108 14736
rect 11868 14714 11892 14716
rect 11948 14714 11972 14716
rect 12028 14714 12052 14716
rect 11890 14662 11892 14714
rect 11954 14662 11966 14714
rect 12028 14662 12030 14714
rect 11868 14660 11892 14662
rect 11948 14660 11972 14662
rect 12028 14660 12052 14662
rect 11812 14640 12108 14660
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 12176 14074 12204 14486
rect 12820 14346 12848 14894
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 12808 14340 12860 14346
rect 12808 14282 12860 14288
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 9784 11886 9996 11914
rect 10704 11898 10732 12786
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 10060 10810 10088 11494
rect 10612 11150 10640 11630
rect 10704 11558 10732 11834
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8864 10266 8892 10474
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8772 8022 8800 8434
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8864 6186 8892 7278
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8680 4690 8708 5782
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8680 4078 8708 4626
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8956 3942 8984 10066
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9098 9820 9394 9840
rect 9154 9818 9178 9820
rect 9234 9818 9258 9820
rect 9314 9818 9338 9820
rect 9176 9766 9178 9818
rect 9240 9766 9252 9818
rect 9314 9766 9316 9818
rect 9154 9764 9178 9766
rect 9234 9764 9258 9766
rect 9314 9764 9338 9766
rect 9098 9744 9394 9764
rect 9098 8732 9394 8752
rect 9154 8730 9178 8732
rect 9234 8730 9258 8732
rect 9314 8730 9338 8732
rect 9176 8678 9178 8730
rect 9240 8678 9252 8730
rect 9314 8678 9316 8730
rect 9154 8676 9178 8678
rect 9234 8676 9258 8678
rect 9314 8676 9338 8678
rect 9098 8656 9394 8676
rect 9508 7954 9536 9930
rect 9692 8634 9720 10542
rect 10060 10538 10088 10746
rect 10612 10538 10640 11086
rect 10704 10606 10732 11494
rect 10796 10996 10824 13126
rect 11348 12782 11376 13670
rect 11812 13628 12108 13648
rect 11868 13626 11892 13628
rect 11948 13626 11972 13628
rect 12028 13626 12052 13628
rect 11890 13574 11892 13626
rect 11954 13574 11966 13626
rect 12028 13574 12030 13626
rect 11868 13572 11892 13574
rect 11948 13572 11972 13574
rect 12028 13572 12052 13574
rect 11812 13552 12108 13572
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 11762 11468 12582
rect 11624 12306 11652 13126
rect 11716 12442 11744 13398
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 11812 12540 12108 12560
rect 11868 12538 11892 12540
rect 11948 12538 11972 12540
rect 12028 12538 12052 12540
rect 11890 12486 11892 12538
rect 11954 12486 11966 12538
rect 12028 12486 12030 12538
rect 11868 12484 11892 12486
rect 11948 12484 11972 12486
rect 12028 12484 12052 12486
rect 11812 12464 12108 12484
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10876 11008 10928 11014
rect 10796 10968 10876 10996
rect 10796 10606 10824 10968
rect 10876 10950 10928 10956
rect 11072 10810 11100 11086
rect 11348 10810 11376 11222
rect 11440 11150 11468 11698
rect 12084 11694 12112 12038
rect 12360 11694 12388 12242
rect 12452 11694 12480 12378
rect 12728 11898 12756 13262
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12084 11540 12112 11630
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 12084 11512 12204 11540
rect 11812 11452 12108 11472
rect 11868 11450 11892 11452
rect 11948 11450 11972 11452
rect 12028 11450 12052 11452
rect 11890 11398 11892 11450
rect 11954 11398 11966 11450
rect 12028 11398 12030 11450
rect 11868 11396 11892 11398
rect 11948 11396 11972 11398
rect 12028 11396 12052 11398
rect 11812 11376 12108 11396
rect 12176 11354 12204 11512
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12268 11218 12296 11562
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11440 10674 11468 11086
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 11716 10266 11744 11086
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10674 12480 10950
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 11812 10364 12108 10384
rect 11868 10362 11892 10364
rect 11948 10362 11972 10364
rect 12028 10362 12052 10364
rect 11890 10310 11892 10362
rect 11954 10310 11966 10362
rect 12028 10310 12030 10362
rect 11868 10308 11892 10310
rect 11948 10308 11972 10310
rect 12028 10308 12052 10310
rect 11812 10288 12108 10308
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 12820 10130 12848 14282
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12912 12442 12940 14214
rect 13004 13394 13032 14826
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13188 14550 13216 14758
rect 13176 14544 13228 14550
rect 13176 14486 13228 14492
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13096 14074 13124 14350
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13280 13734 13308 14010
rect 13372 13802 13400 15506
rect 13832 15094 13860 17711
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14108 16574 14136 17070
rect 14016 16546 14136 16574
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13832 14822 13860 14894
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13924 14618 13952 15982
rect 14016 15502 14044 16546
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 14016 14822 14044 15438
rect 14108 15162 14136 15914
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13372 13394 13400 13738
rect 13648 13530 13676 14214
rect 13924 14074 13952 14554
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13832 13870 13860 13942
rect 14108 13938 14136 15098
rect 14292 15042 14320 15846
rect 14384 15144 14412 18686
rect 14526 18524 14822 18544
rect 14582 18522 14606 18524
rect 14662 18522 14686 18524
rect 14742 18522 14766 18524
rect 14604 18470 14606 18522
rect 14668 18470 14680 18522
rect 14742 18470 14744 18522
rect 14582 18468 14606 18470
rect 14662 18468 14686 18470
rect 14742 18468 14766 18470
rect 14526 18448 14822 18468
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15304 18222 15332 18362
rect 16488 18352 16540 18358
rect 16488 18294 16540 18300
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14526 17436 14822 17456
rect 14582 17434 14606 17436
rect 14662 17434 14686 17436
rect 14742 17434 14766 17436
rect 14604 17382 14606 17434
rect 14668 17382 14680 17434
rect 14742 17382 14744 17434
rect 14582 17380 14606 17382
rect 14662 17380 14686 17382
rect 14742 17380 14766 17382
rect 14526 17360 14822 17380
rect 14936 17202 14964 18022
rect 15120 17882 15148 18158
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15120 17610 15148 17818
rect 15212 17746 15240 18090
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 15304 17082 15332 18158
rect 15396 17542 15424 18158
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15212 17054 15332 17082
rect 15212 16658 15240 17054
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 14526 16348 14822 16368
rect 14582 16346 14606 16348
rect 14662 16346 14686 16348
rect 14742 16346 14766 16348
rect 14604 16294 14606 16346
rect 14668 16294 14680 16346
rect 14742 16294 14744 16346
rect 14582 16292 14606 16294
rect 14662 16292 14686 16294
rect 14742 16292 14766 16294
rect 14526 16272 14822 16292
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 14924 15972 14976 15978
rect 14924 15914 14976 15920
rect 14526 15260 14822 15280
rect 14582 15258 14606 15260
rect 14662 15258 14686 15260
rect 14742 15258 14766 15260
rect 14604 15206 14606 15258
rect 14668 15206 14680 15258
rect 14742 15206 14744 15258
rect 14582 15204 14606 15206
rect 14662 15204 14686 15206
rect 14742 15204 14766 15206
rect 14526 15184 14822 15204
rect 14384 15116 14504 15144
rect 14200 15026 14320 15042
rect 14188 15020 14320 15026
rect 14240 15014 14320 15020
rect 14188 14962 14240 14968
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14384 14074 14412 14826
rect 14476 14482 14504 15116
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14844 14822 14872 14962
rect 14936 14822 14964 15914
rect 15028 15366 15056 15982
rect 15212 15638 15240 16390
rect 15304 16250 15332 16934
rect 15396 16794 15424 17478
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15200 15632 15252 15638
rect 15200 15574 15252 15580
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14936 14482 14964 14758
rect 15028 14618 15056 15302
rect 15488 15026 15516 18022
rect 16500 17882 16528 18294
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15580 17338 15608 17614
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15936 17060 15988 17066
rect 15936 17002 15988 17008
rect 15948 16794 15976 17002
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16132 16522 16160 16594
rect 16120 16516 16172 16522
rect 16120 16458 16172 16464
rect 16132 16046 16160 16458
rect 16592 16114 16620 19892
rect 17972 17746 18000 19892
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16224 15638 16252 15846
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16394 15056 16450 15065
rect 15476 15020 15528 15026
rect 16394 14991 16450 15000
rect 15476 14962 15528 14968
rect 16408 14958 16436 14991
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 15028 14414 15056 14554
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 14526 14172 14822 14192
rect 14582 14170 14606 14172
rect 14662 14170 14686 14172
rect 14742 14170 14766 14172
rect 14604 14118 14606 14170
rect 14668 14118 14680 14170
rect 14742 14118 14744 14170
rect 14582 14116 14606 14118
rect 14662 14116 14686 14118
rect 14742 14116 14766 14118
rect 14526 14096 14822 14116
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13832 13258 13860 13806
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13648 12442 13676 12650
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13832 12102 13860 13194
rect 14526 13084 14822 13104
rect 14582 13082 14606 13084
rect 14662 13082 14686 13084
rect 14742 13082 14766 13084
rect 14604 13030 14606 13082
rect 14668 13030 14680 13082
rect 14742 13030 14744 13082
rect 14582 13028 14606 13030
rect 14662 13028 14686 13030
rect 14742 13028 14766 13030
rect 14526 13008 14822 13028
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 13924 12442 13952 12650
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13372 11218 13400 12038
rect 14526 11996 14822 12016
rect 14582 11994 14606 11996
rect 14662 11994 14686 11996
rect 14742 11994 14766 11996
rect 14604 11942 14606 11994
rect 14668 11942 14680 11994
rect 14742 11942 14744 11994
rect 14582 11940 14606 11942
rect 14662 11940 14686 11942
rect 14742 11940 14766 11942
rect 14526 11920 14822 11940
rect 14936 11762 14964 12650
rect 15120 12345 15148 13806
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15212 12374 15240 13194
rect 15200 12368 15252 12374
rect 15106 12336 15162 12345
rect 15200 12310 15252 12316
rect 15106 12271 15162 12280
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13832 11354 13860 11562
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13096 10538 13124 11018
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9968 9042 9996 9522
rect 10612 9518 10640 9590
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9784 8430 9812 8978
rect 10428 8974 10456 9318
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10428 8634 10456 8910
rect 10520 8634 10548 9386
rect 10612 9178 10640 9454
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 10428 8362 10456 8570
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9968 8022 9996 8230
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 9098 7644 9394 7664
rect 9154 7642 9178 7644
rect 9234 7642 9258 7644
rect 9314 7642 9338 7644
rect 9176 7590 9178 7642
rect 9240 7590 9252 7642
rect 9314 7590 9316 7642
rect 9154 7588 9178 7590
rect 9234 7588 9258 7590
rect 9314 7588 9338 7590
rect 9098 7568 9394 7588
rect 9692 7410 9720 7686
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9098 6556 9394 6576
rect 9154 6554 9178 6556
rect 9234 6554 9258 6556
rect 9314 6554 9338 6556
rect 9176 6502 9178 6554
rect 9240 6502 9252 6554
rect 9314 6502 9316 6554
rect 9154 6500 9178 6502
rect 9234 6500 9258 6502
rect 9314 6500 9338 6502
rect 9098 6480 9394 6500
rect 9508 6338 9536 7142
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9416 6322 9536 6338
rect 9404 6316 9536 6322
rect 9456 6310 9536 6316
rect 9404 6258 9456 6264
rect 9784 6186 9812 6598
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9098 5468 9394 5488
rect 9154 5466 9178 5468
rect 9234 5466 9258 5468
rect 9314 5466 9338 5468
rect 9176 5414 9178 5466
rect 9240 5414 9252 5466
rect 9314 5414 9316 5466
rect 9154 5412 9178 5414
rect 9234 5412 9258 5414
rect 9314 5412 9338 5414
rect 9098 5392 9394 5412
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9508 4826 9536 5034
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9098 4380 9394 4400
rect 9154 4378 9178 4380
rect 9234 4378 9258 4380
rect 9314 4378 9338 4380
rect 9176 4326 9178 4378
rect 9240 4326 9252 4378
rect 9314 4326 9316 4378
rect 9154 4324 9178 4326
rect 9234 4324 9258 4326
rect 9314 4324 9338 4326
rect 9098 4304 9394 4324
rect 9692 4078 9720 4966
rect 9784 4758 9812 5646
rect 10244 5234 10272 6054
rect 10336 5914 10364 7278
rect 10428 6866 10456 7686
rect 10520 7546 10548 8366
rect 10612 8294 10640 8910
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10612 7886 10640 8230
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10796 7546 10824 7958
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 11072 7342 11100 8026
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10612 5778 10640 6666
rect 11164 6458 11192 10066
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 11812 9276 12108 9296
rect 11868 9274 11892 9276
rect 11948 9274 11972 9276
rect 12028 9274 12052 9276
rect 11890 9222 11892 9274
rect 11954 9222 11966 9274
rect 12028 9222 12030 9274
rect 11868 9220 11892 9222
rect 11948 9220 11972 9222
rect 12028 9220 12052 9222
rect 11812 9200 12108 9220
rect 12176 9110 12204 9318
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 11812 8188 12108 8208
rect 11868 8186 11892 8188
rect 11948 8186 11972 8188
rect 12028 8186 12052 8188
rect 11890 8134 11892 8186
rect 11954 8134 11966 8186
rect 12028 8134 12030 8186
rect 11868 8132 11892 8134
rect 11948 8132 11972 8134
rect 12028 8132 12052 8134
rect 11812 8112 12108 8132
rect 12176 8072 12204 8366
rect 12360 8294 12388 9590
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12348 8288 12400 8294
rect 12348 8230 12400 8236
rect 12084 8044 12204 8072
rect 12084 7410 12112 8044
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11812 7100 12108 7120
rect 11868 7098 11892 7100
rect 11948 7098 11972 7100
rect 12028 7098 12052 7100
rect 11890 7046 11892 7098
rect 11954 7046 11966 7098
rect 12028 7046 12030 7098
rect 11868 7044 11892 7046
rect 11948 7044 11972 7046
rect 12028 7044 12052 7046
rect 11812 7024 12108 7044
rect 12176 7002 12204 7686
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12176 6798 12204 6938
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 12268 6662 12296 7754
rect 12360 7342 12388 8230
rect 12452 8022 12480 9454
rect 12820 8974 12848 10066
rect 13188 9178 13216 10066
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13280 9586 13308 9862
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13372 9042 13400 11154
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13648 10062 13676 10678
rect 14016 10606 14044 11494
rect 14936 11218 14964 11698
rect 15212 11286 15240 12310
rect 15200 11280 15252 11286
rect 15200 11222 15252 11228
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 14526 10908 14822 10928
rect 14582 10906 14606 10908
rect 14662 10906 14686 10908
rect 14742 10906 14766 10908
rect 14604 10854 14606 10906
rect 14668 10854 14680 10906
rect 14742 10854 14744 10906
rect 14582 10852 14606 10854
rect 14662 10852 14686 10854
rect 14742 10852 14766 10854
rect 14526 10832 14822 10852
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 14936 10130 14964 10406
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 14526 9820 14822 9840
rect 14582 9818 14606 9820
rect 14662 9818 14686 9820
rect 14742 9818 14766 9820
rect 14604 9766 14606 9818
rect 14668 9766 14680 9818
rect 14742 9766 14744 9818
rect 14582 9764 14606 9766
rect 14662 9764 14686 9766
rect 14742 9764 14766 9766
rect 14526 9744 14822 9764
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13832 9178 13860 9386
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 14936 9042 14964 9318
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12820 8634 12848 8910
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12544 7750 12572 8026
rect 12820 7886 12848 8230
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6866 12480 7142
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 12268 6254 12296 6598
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 11532 5914 11560 6054
rect 11812 6012 12108 6032
rect 11868 6010 11892 6012
rect 11948 6010 11972 6012
rect 12028 6010 12052 6012
rect 11890 5958 11892 6010
rect 11954 5958 11966 6010
rect 12028 5958 12030 6010
rect 11868 5956 11892 5958
rect 11948 5956 11972 5958
rect 12028 5956 12052 5958
rect 11812 5936 12108 5956
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9784 4622 9812 4694
rect 10244 4690 10272 5170
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10520 4758 10548 4966
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9508 3942 9536 4014
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 6012 2650 6040 3334
rect 6384 2748 6680 2768
rect 6440 2746 6464 2748
rect 6520 2746 6544 2748
rect 6600 2746 6624 2748
rect 6462 2694 6464 2746
rect 6526 2694 6538 2746
rect 6600 2694 6602 2746
rect 6440 2692 6464 2694
rect 6520 2692 6544 2694
rect 6600 2692 6624 2694
rect 6384 2672 6680 2692
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 6012 2514 6040 2586
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 7300 898 7328 3334
rect 7392 2650 7420 3470
rect 7760 3194 7788 3470
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 8220 2922 8248 3334
rect 8496 3058 8524 3334
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 8588 2514 8616 3470
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 7300 870 7420 898
rect 7392 800 7420 870
rect 8772 800 8800 3402
rect 9098 3292 9394 3312
rect 9154 3290 9178 3292
rect 9234 3290 9258 3292
rect 9314 3290 9338 3292
rect 9176 3238 9178 3290
rect 9240 3238 9252 3290
rect 9314 3238 9316 3290
rect 9154 3236 9178 3238
rect 9234 3236 9258 3238
rect 9314 3236 9338 3238
rect 9098 3216 9394 3236
rect 9508 3194 9536 3878
rect 9588 3664 9640 3670
rect 9588 3606 9640 3612
rect 9600 3398 9628 3606
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9692 2650 9720 2858
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9784 2514 9812 4558
rect 10612 4078 10640 5510
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 9968 3942 9996 4014
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9968 3738 9996 3878
rect 10612 3738 10640 4014
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 9968 3602 9996 3674
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 10612 2650 10640 2858
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9098 2204 9394 2224
rect 9154 2202 9178 2204
rect 9234 2202 9258 2204
rect 9314 2202 9338 2204
rect 9176 2150 9178 2202
rect 9240 2150 9252 2202
rect 9314 2150 9316 2202
rect 9154 2148 9178 2150
rect 9234 2148 9258 2150
rect 9314 2148 9338 2150
rect 9098 2128 9394 2148
rect 10704 898 10732 5714
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 11072 5370 11100 5578
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11072 5030 11100 5306
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 12072 5228 12124 5234
rect 12176 5216 12204 6054
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12452 5234 12480 5510
rect 12728 5370 12756 5714
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12124 5188 12204 5216
rect 12440 5228 12492 5234
rect 12072 5170 12124 5176
rect 12440 5170 12492 5176
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11072 2582 11100 3334
rect 11256 3058 11284 5170
rect 12820 5114 12848 5714
rect 12636 5098 12848 5114
rect 12624 5092 12848 5098
rect 12676 5086 12848 5092
rect 12624 5034 12676 5040
rect 11812 4924 12108 4944
rect 11868 4922 11892 4924
rect 11948 4922 11972 4924
rect 12028 4922 12052 4924
rect 11890 4870 11892 4922
rect 11954 4870 11966 4922
rect 12028 4870 12030 4922
rect 11868 4868 11892 4870
rect 11948 4868 11972 4870
rect 12028 4868 12052 4870
rect 11812 4848 12108 4868
rect 12820 4826 12848 5086
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12084 4282 12112 4694
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11812 3836 12108 3856
rect 11868 3834 11892 3836
rect 11948 3834 11972 3836
rect 12028 3834 12052 3836
rect 11890 3782 11892 3834
rect 11954 3782 11966 3834
rect 12028 3782 12030 3834
rect 11868 3780 11892 3782
rect 11948 3780 11972 3782
rect 12028 3780 12052 3782
rect 11812 3760 12108 3780
rect 12176 3602 12204 4422
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12544 3670 12572 4082
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 11440 3194 11468 3538
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11440 2650 11468 3130
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11440 2378 11468 2586
rect 11624 2514 11652 3538
rect 11716 3058 11744 3538
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 12176 2854 12204 3538
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 11812 2748 12108 2768
rect 11868 2746 11892 2748
rect 11948 2746 11972 2748
rect 12028 2746 12052 2748
rect 11890 2694 11892 2746
rect 11954 2694 11966 2746
rect 12028 2694 12030 2746
rect 11868 2692 11892 2694
rect 11948 2692 11972 2694
rect 12028 2692 12052 2694
rect 11812 2672 12108 2692
rect 12268 2650 12296 2926
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11428 2372 11480 2378
rect 11428 2314 11480 2320
rect 10612 870 10732 898
rect 10612 800 10640 870
rect 12452 800 12480 3538
rect 12728 2378 12756 3878
rect 13004 3738 13032 8978
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13096 6866 13124 7822
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13188 6254 13216 7958
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13268 7268 13320 7274
rect 13268 7210 13320 7216
rect 13280 7002 13308 7210
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13372 6866 13400 7686
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13556 6730 13584 8434
rect 13740 8022 13768 8910
rect 14526 8732 14822 8752
rect 14582 8730 14606 8732
rect 14662 8730 14686 8732
rect 14742 8730 14766 8732
rect 14604 8678 14606 8730
rect 14668 8678 14680 8730
rect 14742 8678 14744 8730
rect 14582 8676 14606 8678
rect 14662 8676 14686 8678
rect 14742 8676 14766 8678
rect 14526 8656 14822 8676
rect 14936 8498 14964 8978
rect 15212 8634 15240 10950
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15304 9110 15332 9862
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13832 8090 13860 8298
rect 14936 8090 14964 8434
rect 15396 8412 15424 13942
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15948 12306 15976 13126
rect 16040 12782 16068 13670
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15488 10810 15516 11562
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15488 9586 15516 10066
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15580 9518 15608 10066
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15764 8566 15792 10134
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15856 9722 15884 10066
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15856 8634 15884 9658
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15948 9178 15976 9454
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15476 8560 15528 8566
rect 15752 8560 15804 8566
rect 15476 8502 15528 8508
rect 15672 8508 15752 8514
rect 15672 8502 15804 8508
rect 15212 8384 15424 8412
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 14526 7644 14822 7664
rect 14582 7642 14606 7644
rect 14662 7642 14686 7644
rect 14742 7642 14766 7644
rect 14604 7590 14606 7642
rect 14668 7590 14680 7642
rect 14742 7590 14744 7642
rect 14582 7588 14606 7590
rect 14662 7588 14686 7590
rect 14742 7588 14766 7590
rect 14526 7568 14822 7588
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13544 6724 13596 6730
rect 13544 6666 13596 6672
rect 13832 6458 13860 7210
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14384 6254 14412 6666
rect 14526 6556 14822 6576
rect 14582 6554 14606 6556
rect 14662 6554 14686 6556
rect 14742 6554 14766 6556
rect 14604 6502 14606 6554
rect 14668 6502 14680 6554
rect 14742 6502 14744 6554
rect 14582 6500 14606 6502
rect 14662 6500 14686 6502
rect 14742 6500 14766 6502
rect 14526 6480 14822 6500
rect 14936 6458 14964 6802
rect 15028 6458 15056 7142
rect 15212 6746 15240 8384
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15120 6718 15240 6746
rect 15120 6662 15148 6718
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 15028 6118 15056 6394
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 14108 5710 14136 6054
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14108 5234 14136 5646
rect 14384 5370 14412 6054
rect 15212 5846 15240 6598
rect 15304 5914 15332 7890
rect 15488 7818 15516 8502
rect 15672 8486 15792 8502
rect 15568 8424 15620 8430
rect 15672 8412 15700 8486
rect 15620 8384 15700 8412
rect 15568 8366 15620 8372
rect 15672 8090 15700 8384
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15476 7812 15528 7818
rect 15476 7754 15528 7760
rect 15856 7342 15884 8230
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15396 6254 15424 6802
rect 15580 6458 15608 6802
rect 15948 6798 15976 7278
rect 16132 6866 16160 14758
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16224 12374 16252 14214
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16316 13258 16344 13806
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 16316 11676 16344 13194
rect 16408 12986 16436 13330
rect 16500 13190 16528 13466
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16408 12442 16436 12922
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16500 12306 16528 13126
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16592 12442 16620 12786
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 16396 11688 16448 11694
rect 16316 11648 16396 11676
rect 16396 11630 16448 11636
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 11286 16252 11494
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16408 10130 16436 11630
rect 16500 11354 16528 12242
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 9042 16344 9862
rect 16394 9616 16450 9625
rect 16394 9551 16450 9560
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16408 8430 16436 9551
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16684 7585 16712 7890
rect 16670 7576 16726 7585
rect 16670 7511 16726 7520
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15580 5914 15608 6190
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15200 5840 15252 5846
rect 15672 5794 15700 6734
rect 16224 6458 16252 7346
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 15200 5782 15252 5788
rect 15580 5766 15700 5794
rect 16212 5840 16264 5846
rect 16212 5782 16264 5788
rect 14526 5468 14822 5488
rect 14582 5466 14606 5468
rect 14662 5466 14686 5468
rect 14742 5466 14766 5468
rect 14604 5414 14606 5466
rect 14668 5414 14680 5466
rect 14742 5414 14744 5466
rect 14582 5412 14606 5414
rect 14662 5412 14686 5414
rect 14742 5412 14766 5414
rect 14526 5392 14822 5412
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 13360 5092 13412 5098
rect 13360 5034 13412 5040
rect 13372 4826 13400 5034
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13360 4684 13412 4690
rect 13360 4626 13412 4632
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 13372 3670 13400 4626
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13740 3738 13768 3946
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 13372 2990 13400 3606
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13188 2582 13216 2790
rect 13740 2582 13768 3402
rect 13832 3194 13860 4558
rect 14108 4146 14136 5170
rect 15016 5092 15068 5098
rect 15016 5034 15068 5040
rect 15028 4826 15056 5034
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 14526 4380 14822 4400
rect 14582 4378 14606 4380
rect 14662 4378 14686 4380
rect 14742 4378 14766 4380
rect 14604 4326 14606 4378
rect 14668 4326 14680 4378
rect 14742 4326 14744 4378
rect 14582 4324 14606 4326
rect 14662 4324 14686 4326
rect 14742 4324 14766 4326
rect 14526 4304 14822 4324
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 14108 2514 14136 4082
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 14200 3194 14228 3946
rect 14936 3602 14964 4082
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14526 3292 14822 3312
rect 14582 3290 14606 3292
rect 14662 3290 14686 3292
rect 14742 3290 14766 3292
rect 14604 3238 14606 3290
rect 14668 3238 14680 3290
rect 14742 3238 14744 3290
rect 14582 3236 14606 3238
rect 14662 3236 14686 3238
rect 14742 3236 14766 3238
rect 14526 3216 14822 3236
rect 15028 3194 15056 3878
rect 15212 3670 15240 4626
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15304 3942 15332 4218
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15212 3194 15240 3470
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 15016 3188 15068 3194
rect 15016 3130 15068 3136
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15028 3058 15056 3130
rect 15580 3126 15608 5766
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 12716 2372 12768 2378
rect 12716 2314 12768 2320
rect 14292 800 14320 2926
rect 15028 2854 15056 2994
rect 15476 2916 15528 2922
rect 15476 2858 15528 2864
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15488 2650 15516 2858
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15580 2582 15608 3062
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 15672 2514 15700 4422
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 14526 2204 14822 2224
rect 14582 2202 14606 2204
rect 14662 2202 14686 2204
rect 14742 2202 14766 2204
rect 14604 2150 14606 2202
rect 14668 2150 14680 2202
rect 14742 2150 14744 2202
rect 14582 2148 14606 2150
rect 14662 2148 14686 2150
rect 14742 2148 14766 2150
rect 14526 2128 14822 2148
rect 15764 2145 15792 4626
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15856 3534 15884 4014
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15856 2990 15884 3470
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15948 2774 15976 5510
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 16040 4282 16068 4966
rect 16224 4826 16252 5782
rect 16408 4865 16436 6190
rect 16394 4856 16450 4865
rect 16212 4820 16264 4826
rect 16394 4791 16450 4800
rect 16212 4762 16264 4768
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 16040 2990 16068 4218
rect 16408 4078 16436 4626
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 16224 3670 16252 3878
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 15948 2746 16160 2774
rect 15750 2136 15806 2145
rect 15750 2071 15806 2080
rect 16132 800 16160 2746
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16500 2106 16528 2246
rect 16488 2100 16540 2106
rect 16488 2042 16540 2048
rect 17512 800 17540 2450
rect 478 0 534 800
rect 1858 0 1914 800
rect 3698 0 3754 800
rect 5538 0 5594 800
rect 7378 0 7434 800
rect 8758 0 8814 800
rect 10598 0 10654 800
rect 12438 0 12494 800
rect 14278 0 14334 800
rect 16118 0 16174 800
rect 17498 0 17554 800
<< via2 >>
rect 1766 18400 1822 18456
rect 3670 18522 3726 18524
rect 3750 18522 3806 18524
rect 3830 18522 3886 18524
rect 3910 18522 3966 18524
rect 3670 18470 3696 18522
rect 3696 18470 3726 18522
rect 3750 18470 3760 18522
rect 3760 18470 3806 18522
rect 3830 18470 3876 18522
rect 3876 18470 3886 18522
rect 3910 18470 3940 18522
rect 3940 18470 3966 18522
rect 3670 18468 3726 18470
rect 3750 18468 3806 18470
rect 3830 18468 3886 18470
rect 3910 18468 3966 18470
rect 1950 15680 2006 15736
rect 2778 12960 2834 13016
rect 1766 10920 1822 10976
rect 1950 8200 2006 8256
rect 3670 17434 3726 17436
rect 3750 17434 3806 17436
rect 3830 17434 3886 17436
rect 3910 17434 3966 17436
rect 3670 17382 3696 17434
rect 3696 17382 3726 17434
rect 3750 17382 3760 17434
rect 3760 17382 3806 17434
rect 3830 17382 3876 17434
rect 3876 17382 3886 17434
rect 3910 17382 3940 17434
rect 3940 17382 3966 17434
rect 3670 17380 3726 17382
rect 3750 17380 3806 17382
rect 3830 17380 3886 17382
rect 3910 17380 3966 17382
rect 3670 16346 3726 16348
rect 3750 16346 3806 16348
rect 3830 16346 3886 16348
rect 3910 16346 3966 16348
rect 3670 16294 3696 16346
rect 3696 16294 3726 16346
rect 3750 16294 3760 16346
rect 3760 16294 3806 16346
rect 3830 16294 3876 16346
rect 3876 16294 3886 16346
rect 3910 16294 3940 16346
rect 3940 16294 3966 16346
rect 3670 16292 3726 16294
rect 3750 16292 3806 16294
rect 3830 16292 3886 16294
rect 3910 16292 3966 16294
rect 3670 15258 3726 15260
rect 3750 15258 3806 15260
rect 3830 15258 3886 15260
rect 3910 15258 3966 15260
rect 3670 15206 3696 15258
rect 3696 15206 3726 15258
rect 3750 15206 3760 15258
rect 3760 15206 3806 15258
rect 3830 15206 3876 15258
rect 3876 15206 3886 15258
rect 3910 15206 3940 15258
rect 3940 15206 3966 15258
rect 3670 15204 3726 15206
rect 3750 15204 3806 15206
rect 3830 15204 3886 15206
rect 3910 15204 3966 15206
rect 3670 14170 3726 14172
rect 3750 14170 3806 14172
rect 3830 14170 3886 14172
rect 3910 14170 3966 14172
rect 3670 14118 3696 14170
rect 3696 14118 3726 14170
rect 3750 14118 3760 14170
rect 3760 14118 3806 14170
rect 3830 14118 3876 14170
rect 3876 14118 3886 14170
rect 3910 14118 3940 14170
rect 3940 14118 3966 14170
rect 3670 14116 3726 14118
rect 3750 14116 3806 14118
rect 3830 14116 3886 14118
rect 3910 14116 3966 14118
rect 3670 13082 3726 13084
rect 3750 13082 3806 13084
rect 3830 13082 3886 13084
rect 3910 13082 3966 13084
rect 3670 13030 3696 13082
rect 3696 13030 3726 13082
rect 3750 13030 3760 13082
rect 3760 13030 3806 13082
rect 3830 13030 3876 13082
rect 3876 13030 3886 13082
rect 3910 13030 3940 13082
rect 3940 13030 3966 13082
rect 3670 13028 3726 13030
rect 3750 13028 3806 13030
rect 3830 13028 3886 13030
rect 3910 13028 3966 13030
rect 3670 11994 3726 11996
rect 3750 11994 3806 11996
rect 3830 11994 3886 11996
rect 3910 11994 3966 11996
rect 3670 11942 3696 11994
rect 3696 11942 3726 11994
rect 3750 11942 3760 11994
rect 3760 11942 3806 11994
rect 3830 11942 3876 11994
rect 3876 11942 3886 11994
rect 3910 11942 3940 11994
rect 3940 11942 3966 11994
rect 3670 11940 3726 11942
rect 3750 11940 3806 11942
rect 3830 11940 3886 11942
rect 3910 11940 3966 11942
rect 3670 10906 3726 10908
rect 3750 10906 3806 10908
rect 3830 10906 3886 10908
rect 3910 10906 3966 10908
rect 3670 10854 3696 10906
rect 3696 10854 3726 10906
rect 3750 10854 3760 10906
rect 3760 10854 3806 10906
rect 3830 10854 3876 10906
rect 3876 10854 3886 10906
rect 3910 10854 3940 10906
rect 3940 10854 3966 10906
rect 3670 10852 3726 10854
rect 3750 10852 3806 10854
rect 3830 10852 3886 10854
rect 3910 10852 3966 10854
rect 3670 9818 3726 9820
rect 3750 9818 3806 9820
rect 3830 9818 3886 9820
rect 3910 9818 3966 9820
rect 3670 9766 3696 9818
rect 3696 9766 3726 9818
rect 3750 9766 3760 9818
rect 3760 9766 3806 9818
rect 3830 9766 3876 9818
rect 3876 9766 3886 9818
rect 3910 9766 3940 9818
rect 3940 9766 3966 9818
rect 3670 9764 3726 9766
rect 3750 9764 3806 9766
rect 3830 9764 3886 9766
rect 3910 9764 3966 9766
rect 3670 8730 3726 8732
rect 3750 8730 3806 8732
rect 3830 8730 3886 8732
rect 3910 8730 3966 8732
rect 3670 8678 3696 8730
rect 3696 8678 3726 8730
rect 3750 8678 3760 8730
rect 3760 8678 3806 8730
rect 3830 8678 3876 8730
rect 3876 8678 3886 8730
rect 3910 8678 3940 8730
rect 3940 8678 3966 8730
rect 3670 8676 3726 8678
rect 3750 8676 3806 8678
rect 3830 8676 3886 8678
rect 3910 8676 3966 8678
rect 3670 7642 3726 7644
rect 3750 7642 3806 7644
rect 3830 7642 3886 7644
rect 3910 7642 3966 7644
rect 3670 7590 3696 7642
rect 3696 7590 3726 7642
rect 3750 7590 3760 7642
rect 3760 7590 3806 7642
rect 3830 7590 3876 7642
rect 3876 7590 3886 7642
rect 3910 7590 3940 7642
rect 3940 7590 3966 7642
rect 3670 7588 3726 7590
rect 3750 7588 3806 7590
rect 3830 7588 3886 7590
rect 3910 7588 3966 7590
rect 1398 5480 1454 5536
rect 3670 6554 3726 6556
rect 3750 6554 3806 6556
rect 3830 6554 3886 6556
rect 3910 6554 3966 6556
rect 3670 6502 3696 6554
rect 3696 6502 3726 6554
rect 3750 6502 3760 6554
rect 3760 6502 3806 6554
rect 3830 6502 3876 6554
rect 3876 6502 3886 6554
rect 3910 6502 3940 6554
rect 3940 6502 3966 6554
rect 3670 6500 3726 6502
rect 3750 6500 3806 6502
rect 3830 6500 3886 6502
rect 3910 6500 3966 6502
rect 3670 5466 3726 5468
rect 3750 5466 3806 5468
rect 3830 5466 3886 5468
rect 3910 5466 3966 5468
rect 3670 5414 3696 5466
rect 3696 5414 3726 5466
rect 3750 5414 3760 5466
rect 3760 5414 3806 5466
rect 3830 5414 3876 5466
rect 3876 5414 3886 5466
rect 3910 5414 3940 5466
rect 3940 5414 3966 5466
rect 3670 5412 3726 5414
rect 3750 5412 3806 5414
rect 3830 5412 3886 5414
rect 3910 5412 3966 5414
rect 3670 4378 3726 4380
rect 3750 4378 3806 4380
rect 3830 4378 3886 4380
rect 3910 4378 3966 4380
rect 3670 4326 3696 4378
rect 3696 4326 3726 4378
rect 3750 4326 3760 4378
rect 3760 4326 3806 4378
rect 3830 4326 3876 4378
rect 3876 4326 3886 4378
rect 3910 4326 3940 4378
rect 3940 4326 3966 4378
rect 3670 4324 3726 4326
rect 3750 4324 3806 4326
rect 3830 4324 3886 4326
rect 3910 4324 3966 4326
rect 3670 3290 3726 3292
rect 3750 3290 3806 3292
rect 3830 3290 3886 3292
rect 3910 3290 3966 3292
rect 3670 3238 3696 3290
rect 3696 3238 3726 3290
rect 3750 3238 3760 3290
rect 3760 3238 3806 3290
rect 3830 3238 3876 3290
rect 3876 3238 3886 3290
rect 3910 3238 3940 3290
rect 3940 3238 3966 3290
rect 3670 3236 3726 3238
rect 3750 3236 3806 3238
rect 3830 3236 3886 3238
rect 3910 3236 3966 3238
rect 3974 2760 4030 2816
rect 3670 2202 3726 2204
rect 3750 2202 3806 2204
rect 3830 2202 3886 2204
rect 3910 2202 3966 2204
rect 3670 2150 3696 2202
rect 3696 2150 3726 2202
rect 3750 2150 3760 2202
rect 3760 2150 3806 2202
rect 3830 2150 3876 2202
rect 3876 2150 3886 2202
rect 3910 2150 3940 2202
rect 3940 2150 3966 2202
rect 3670 2148 3726 2150
rect 3750 2148 3806 2150
rect 3830 2148 3886 2150
rect 3910 2148 3966 2150
rect 9098 18522 9154 18524
rect 9178 18522 9234 18524
rect 9258 18522 9314 18524
rect 9338 18522 9394 18524
rect 9098 18470 9124 18522
rect 9124 18470 9154 18522
rect 9178 18470 9188 18522
rect 9188 18470 9234 18522
rect 9258 18470 9304 18522
rect 9304 18470 9314 18522
rect 9338 18470 9368 18522
rect 9368 18470 9394 18522
rect 9098 18468 9154 18470
rect 9178 18468 9234 18470
rect 9258 18468 9314 18470
rect 9338 18468 9394 18470
rect 6384 17978 6440 17980
rect 6464 17978 6520 17980
rect 6544 17978 6600 17980
rect 6624 17978 6680 17980
rect 6384 17926 6410 17978
rect 6410 17926 6440 17978
rect 6464 17926 6474 17978
rect 6474 17926 6520 17978
rect 6544 17926 6590 17978
rect 6590 17926 6600 17978
rect 6624 17926 6654 17978
rect 6654 17926 6680 17978
rect 6384 17924 6440 17926
rect 6464 17924 6520 17926
rect 6544 17924 6600 17926
rect 6624 17924 6680 17926
rect 6384 16890 6440 16892
rect 6464 16890 6520 16892
rect 6544 16890 6600 16892
rect 6624 16890 6680 16892
rect 6384 16838 6410 16890
rect 6410 16838 6440 16890
rect 6464 16838 6474 16890
rect 6474 16838 6520 16890
rect 6544 16838 6590 16890
rect 6590 16838 6600 16890
rect 6624 16838 6654 16890
rect 6654 16838 6680 16890
rect 6384 16836 6440 16838
rect 6464 16836 6520 16838
rect 6544 16836 6600 16838
rect 6624 16836 6680 16838
rect 6384 15802 6440 15804
rect 6464 15802 6520 15804
rect 6544 15802 6600 15804
rect 6624 15802 6680 15804
rect 6384 15750 6410 15802
rect 6410 15750 6440 15802
rect 6464 15750 6474 15802
rect 6474 15750 6520 15802
rect 6544 15750 6590 15802
rect 6590 15750 6600 15802
rect 6624 15750 6654 15802
rect 6654 15750 6680 15802
rect 6384 15748 6440 15750
rect 6464 15748 6520 15750
rect 6544 15748 6600 15750
rect 6624 15748 6680 15750
rect 6384 14714 6440 14716
rect 6464 14714 6520 14716
rect 6544 14714 6600 14716
rect 6624 14714 6680 14716
rect 6384 14662 6410 14714
rect 6410 14662 6440 14714
rect 6464 14662 6474 14714
rect 6474 14662 6520 14714
rect 6544 14662 6590 14714
rect 6590 14662 6600 14714
rect 6624 14662 6654 14714
rect 6654 14662 6680 14714
rect 6384 14660 6440 14662
rect 6464 14660 6520 14662
rect 6544 14660 6600 14662
rect 6624 14660 6680 14662
rect 6384 13626 6440 13628
rect 6464 13626 6520 13628
rect 6544 13626 6600 13628
rect 6624 13626 6680 13628
rect 6384 13574 6410 13626
rect 6410 13574 6440 13626
rect 6464 13574 6474 13626
rect 6474 13574 6520 13626
rect 6544 13574 6590 13626
rect 6590 13574 6600 13626
rect 6624 13574 6654 13626
rect 6654 13574 6680 13626
rect 6384 13572 6440 13574
rect 6464 13572 6520 13574
rect 6544 13572 6600 13574
rect 6624 13572 6680 13574
rect 6384 12538 6440 12540
rect 6464 12538 6520 12540
rect 6544 12538 6600 12540
rect 6624 12538 6680 12540
rect 6384 12486 6410 12538
rect 6410 12486 6440 12538
rect 6464 12486 6474 12538
rect 6474 12486 6520 12538
rect 6544 12486 6590 12538
rect 6590 12486 6600 12538
rect 6624 12486 6654 12538
rect 6654 12486 6680 12538
rect 6384 12484 6440 12486
rect 6464 12484 6520 12486
rect 6544 12484 6600 12486
rect 6624 12484 6680 12486
rect 6384 11450 6440 11452
rect 6464 11450 6520 11452
rect 6544 11450 6600 11452
rect 6624 11450 6680 11452
rect 6384 11398 6410 11450
rect 6410 11398 6440 11450
rect 6464 11398 6474 11450
rect 6474 11398 6520 11450
rect 6544 11398 6590 11450
rect 6590 11398 6600 11450
rect 6624 11398 6654 11450
rect 6654 11398 6680 11450
rect 6384 11396 6440 11398
rect 6464 11396 6520 11398
rect 6544 11396 6600 11398
rect 6624 11396 6680 11398
rect 4710 9560 4766 9616
rect 6384 10362 6440 10364
rect 6464 10362 6520 10364
rect 6544 10362 6600 10364
rect 6624 10362 6680 10364
rect 6384 10310 6410 10362
rect 6410 10310 6440 10362
rect 6464 10310 6474 10362
rect 6474 10310 6520 10362
rect 6544 10310 6590 10362
rect 6590 10310 6600 10362
rect 6624 10310 6654 10362
rect 6654 10310 6680 10362
rect 6384 10308 6440 10310
rect 6464 10308 6520 10310
rect 6544 10308 6600 10310
rect 6624 10308 6680 10310
rect 9098 17434 9154 17436
rect 9178 17434 9234 17436
rect 9258 17434 9314 17436
rect 9338 17434 9394 17436
rect 9098 17382 9124 17434
rect 9124 17382 9154 17434
rect 9178 17382 9188 17434
rect 9188 17382 9234 17434
rect 9258 17382 9304 17434
rect 9304 17382 9314 17434
rect 9338 17382 9368 17434
rect 9368 17382 9394 17434
rect 9098 17380 9154 17382
rect 9178 17380 9234 17382
rect 9258 17380 9314 17382
rect 9338 17380 9394 17382
rect 9098 16346 9154 16348
rect 9178 16346 9234 16348
rect 9258 16346 9314 16348
rect 9338 16346 9394 16348
rect 9098 16294 9124 16346
rect 9124 16294 9154 16346
rect 9178 16294 9188 16346
rect 9188 16294 9234 16346
rect 9258 16294 9304 16346
rect 9304 16294 9314 16346
rect 9338 16294 9368 16346
rect 9368 16294 9394 16346
rect 9098 16292 9154 16294
rect 9178 16292 9234 16294
rect 9258 16292 9314 16294
rect 9338 16292 9394 16294
rect 9098 15258 9154 15260
rect 9178 15258 9234 15260
rect 9258 15258 9314 15260
rect 9338 15258 9394 15260
rect 9098 15206 9124 15258
rect 9124 15206 9154 15258
rect 9178 15206 9188 15258
rect 9188 15206 9234 15258
rect 9258 15206 9304 15258
rect 9304 15206 9314 15258
rect 9338 15206 9368 15258
rect 9368 15206 9394 15258
rect 9098 15204 9154 15206
rect 9178 15204 9234 15206
rect 9258 15204 9314 15206
rect 9338 15204 9394 15206
rect 6384 9274 6440 9276
rect 6464 9274 6520 9276
rect 6544 9274 6600 9276
rect 6624 9274 6680 9276
rect 6384 9222 6410 9274
rect 6410 9222 6440 9274
rect 6464 9222 6474 9274
rect 6474 9222 6520 9274
rect 6544 9222 6590 9274
rect 6590 9222 6600 9274
rect 6624 9222 6654 9274
rect 6654 9222 6680 9274
rect 6384 9220 6440 9222
rect 6464 9220 6520 9222
rect 6544 9220 6600 9222
rect 6624 9220 6680 9222
rect 6384 8186 6440 8188
rect 6464 8186 6520 8188
rect 6544 8186 6600 8188
rect 6624 8186 6680 8188
rect 6384 8134 6410 8186
rect 6410 8134 6440 8186
rect 6464 8134 6474 8186
rect 6474 8134 6520 8186
rect 6544 8134 6590 8186
rect 6590 8134 6600 8186
rect 6624 8134 6654 8186
rect 6654 8134 6680 8186
rect 6384 8132 6440 8134
rect 6464 8132 6520 8134
rect 6544 8132 6600 8134
rect 6624 8132 6680 8134
rect 6384 7098 6440 7100
rect 6464 7098 6520 7100
rect 6544 7098 6600 7100
rect 6624 7098 6680 7100
rect 6384 7046 6410 7098
rect 6410 7046 6440 7098
rect 6464 7046 6474 7098
rect 6474 7046 6520 7098
rect 6544 7046 6590 7098
rect 6590 7046 6600 7098
rect 6624 7046 6654 7098
rect 6654 7046 6680 7098
rect 6384 7044 6440 7046
rect 6464 7044 6520 7046
rect 6544 7044 6600 7046
rect 6624 7044 6680 7046
rect 9098 14170 9154 14172
rect 9178 14170 9234 14172
rect 9258 14170 9314 14172
rect 9338 14170 9394 14172
rect 9098 14118 9124 14170
rect 9124 14118 9154 14170
rect 9178 14118 9188 14170
rect 9188 14118 9234 14170
rect 9258 14118 9304 14170
rect 9304 14118 9314 14170
rect 9338 14118 9368 14170
rect 9368 14118 9394 14170
rect 9098 14116 9154 14118
rect 9178 14116 9234 14118
rect 9258 14116 9314 14118
rect 9338 14116 9394 14118
rect 11812 17978 11868 17980
rect 11892 17978 11948 17980
rect 11972 17978 12028 17980
rect 12052 17978 12108 17980
rect 11812 17926 11838 17978
rect 11838 17926 11868 17978
rect 11892 17926 11902 17978
rect 11902 17926 11948 17978
rect 11972 17926 12018 17978
rect 12018 17926 12028 17978
rect 12052 17926 12082 17978
rect 12082 17926 12108 17978
rect 11812 17924 11868 17926
rect 11892 17924 11948 17926
rect 11972 17924 12028 17926
rect 12052 17924 12108 17926
rect 11812 16890 11868 16892
rect 11892 16890 11948 16892
rect 11972 16890 12028 16892
rect 12052 16890 12108 16892
rect 11812 16838 11838 16890
rect 11838 16838 11868 16890
rect 11892 16838 11902 16890
rect 11902 16838 11948 16890
rect 11972 16838 12018 16890
rect 12018 16838 12028 16890
rect 12052 16838 12082 16890
rect 12082 16838 12108 16890
rect 11812 16836 11868 16838
rect 11892 16836 11948 16838
rect 11972 16836 12028 16838
rect 12052 16836 12108 16838
rect 13818 17720 13874 17776
rect 11812 15802 11868 15804
rect 11892 15802 11948 15804
rect 11972 15802 12028 15804
rect 12052 15802 12108 15804
rect 11812 15750 11838 15802
rect 11838 15750 11868 15802
rect 11892 15750 11902 15802
rect 11902 15750 11948 15802
rect 11972 15750 12018 15802
rect 12018 15750 12028 15802
rect 12052 15750 12082 15802
rect 12082 15750 12108 15802
rect 11812 15748 11868 15750
rect 11892 15748 11948 15750
rect 11972 15748 12028 15750
rect 12052 15748 12108 15750
rect 9098 13082 9154 13084
rect 9178 13082 9234 13084
rect 9258 13082 9314 13084
rect 9338 13082 9394 13084
rect 9098 13030 9124 13082
rect 9124 13030 9154 13082
rect 9178 13030 9188 13082
rect 9188 13030 9234 13082
rect 9258 13030 9304 13082
rect 9304 13030 9314 13082
rect 9338 13030 9368 13082
rect 9368 13030 9394 13082
rect 9098 13028 9154 13030
rect 9178 13028 9234 13030
rect 9258 13028 9314 13030
rect 9338 13028 9394 13030
rect 8574 9560 8630 9616
rect 6384 6010 6440 6012
rect 6464 6010 6520 6012
rect 6544 6010 6600 6012
rect 6624 6010 6680 6012
rect 6384 5958 6410 6010
rect 6410 5958 6440 6010
rect 6464 5958 6474 6010
rect 6474 5958 6520 6010
rect 6544 5958 6590 6010
rect 6590 5958 6600 6010
rect 6624 5958 6654 6010
rect 6654 5958 6680 6010
rect 6384 5956 6440 5958
rect 6464 5956 6520 5958
rect 6544 5956 6600 5958
rect 6624 5956 6680 5958
rect 6384 4922 6440 4924
rect 6464 4922 6520 4924
rect 6544 4922 6600 4924
rect 6624 4922 6680 4924
rect 6384 4870 6410 4922
rect 6410 4870 6440 4922
rect 6464 4870 6474 4922
rect 6474 4870 6520 4922
rect 6544 4870 6590 4922
rect 6590 4870 6600 4922
rect 6624 4870 6654 4922
rect 6654 4870 6680 4922
rect 6384 4868 6440 4870
rect 6464 4868 6520 4870
rect 6544 4868 6600 4870
rect 6624 4868 6680 4870
rect 6384 3834 6440 3836
rect 6464 3834 6520 3836
rect 6544 3834 6600 3836
rect 6624 3834 6680 3836
rect 6384 3782 6410 3834
rect 6410 3782 6440 3834
rect 6464 3782 6474 3834
rect 6474 3782 6520 3834
rect 6544 3782 6590 3834
rect 6590 3782 6600 3834
rect 6624 3782 6654 3834
rect 6654 3782 6680 3834
rect 6384 3780 6440 3782
rect 6464 3780 6520 3782
rect 6544 3780 6600 3782
rect 6624 3780 6680 3782
rect 9098 11994 9154 11996
rect 9178 11994 9234 11996
rect 9258 11994 9314 11996
rect 9338 11994 9394 11996
rect 9098 11942 9124 11994
rect 9124 11942 9154 11994
rect 9178 11942 9188 11994
rect 9188 11942 9234 11994
rect 9258 11942 9304 11994
rect 9304 11942 9314 11994
rect 9338 11942 9368 11994
rect 9368 11942 9394 11994
rect 9098 11940 9154 11942
rect 9178 11940 9234 11942
rect 9258 11940 9314 11942
rect 9338 11940 9394 11942
rect 9098 10906 9154 10908
rect 9178 10906 9234 10908
rect 9258 10906 9314 10908
rect 9338 10906 9394 10908
rect 9098 10854 9124 10906
rect 9124 10854 9154 10906
rect 9178 10854 9188 10906
rect 9188 10854 9234 10906
rect 9258 10854 9304 10906
rect 9304 10854 9314 10906
rect 9338 10854 9368 10906
rect 9368 10854 9394 10906
rect 9098 10852 9154 10854
rect 9178 10852 9234 10854
rect 9258 10852 9314 10854
rect 9338 10852 9394 10854
rect 11812 14714 11868 14716
rect 11892 14714 11948 14716
rect 11972 14714 12028 14716
rect 12052 14714 12108 14716
rect 11812 14662 11838 14714
rect 11838 14662 11868 14714
rect 11892 14662 11902 14714
rect 11902 14662 11948 14714
rect 11972 14662 12018 14714
rect 12018 14662 12028 14714
rect 12052 14662 12082 14714
rect 12082 14662 12108 14714
rect 11812 14660 11868 14662
rect 11892 14660 11948 14662
rect 11972 14660 12028 14662
rect 12052 14660 12108 14662
rect 9098 9818 9154 9820
rect 9178 9818 9234 9820
rect 9258 9818 9314 9820
rect 9338 9818 9394 9820
rect 9098 9766 9124 9818
rect 9124 9766 9154 9818
rect 9178 9766 9188 9818
rect 9188 9766 9234 9818
rect 9258 9766 9304 9818
rect 9304 9766 9314 9818
rect 9338 9766 9368 9818
rect 9368 9766 9394 9818
rect 9098 9764 9154 9766
rect 9178 9764 9234 9766
rect 9258 9764 9314 9766
rect 9338 9764 9394 9766
rect 9098 8730 9154 8732
rect 9178 8730 9234 8732
rect 9258 8730 9314 8732
rect 9338 8730 9394 8732
rect 9098 8678 9124 8730
rect 9124 8678 9154 8730
rect 9178 8678 9188 8730
rect 9188 8678 9234 8730
rect 9258 8678 9304 8730
rect 9304 8678 9314 8730
rect 9338 8678 9368 8730
rect 9368 8678 9394 8730
rect 9098 8676 9154 8678
rect 9178 8676 9234 8678
rect 9258 8676 9314 8678
rect 9338 8676 9394 8678
rect 11812 13626 11868 13628
rect 11892 13626 11948 13628
rect 11972 13626 12028 13628
rect 12052 13626 12108 13628
rect 11812 13574 11838 13626
rect 11838 13574 11868 13626
rect 11892 13574 11902 13626
rect 11902 13574 11948 13626
rect 11972 13574 12018 13626
rect 12018 13574 12028 13626
rect 12052 13574 12082 13626
rect 12082 13574 12108 13626
rect 11812 13572 11868 13574
rect 11892 13572 11948 13574
rect 11972 13572 12028 13574
rect 12052 13572 12108 13574
rect 11812 12538 11868 12540
rect 11892 12538 11948 12540
rect 11972 12538 12028 12540
rect 12052 12538 12108 12540
rect 11812 12486 11838 12538
rect 11838 12486 11868 12538
rect 11892 12486 11902 12538
rect 11902 12486 11948 12538
rect 11972 12486 12018 12538
rect 12018 12486 12028 12538
rect 12052 12486 12082 12538
rect 12082 12486 12108 12538
rect 11812 12484 11868 12486
rect 11892 12484 11948 12486
rect 11972 12484 12028 12486
rect 12052 12484 12108 12486
rect 11812 11450 11868 11452
rect 11892 11450 11948 11452
rect 11972 11450 12028 11452
rect 12052 11450 12108 11452
rect 11812 11398 11838 11450
rect 11838 11398 11868 11450
rect 11892 11398 11902 11450
rect 11902 11398 11948 11450
rect 11972 11398 12018 11450
rect 12018 11398 12028 11450
rect 12052 11398 12082 11450
rect 12082 11398 12108 11450
rect 11812 11396 11868 11398
rect 11892 11396 11948 11398
rect 11972 11396 12028 11398
rect 12052 11396 12108 11398
rect 11812 10362 11868 10364
rect 11892 10362 11948 10364
rect 11972 10362 12028 10364
rect 12052 10362 12108 10364
rect 11812 10310 11838 10362
rect 11838 10310 11868 10362
rect 11892 10310 11902 10362
rect 11902 10310 11948 10362
rect 11972 10310 12018 10362
rect 12018 10310 12028 10362
rect 12052 10310 12082 10362
rect 12082 10310 12108 10362
rect 11812 10308 11868 10310
rect 11892 10308 11948 10310
rect 11972 10308 12028 10310
rect 12052 10308 12108 10310
rect 14526 18522 14582 18524
rect 14606 18522 14662 18524
rect 14686 18522 14742 18524
rect 14766 18522 14822 18524
rect 14526 18470 14552 18522
rect 14552 18470 14582 18522
rect 14606 18470 14616 18522
rect 14616 18470 14662 18522
rect 14686 18470 14732 18522
rect 14732 18470 14742 18522
rect 14766 18470 14796 18522
rect 14796 18470 14822 18522
rect 14526 18468 14582 18470
rect 14606 18468 14662 18470
rect 14686 18468 14742 18470
rect 14766 18468 14822 18470
rect 14526 17434 14582 17436
rect 14606 17434 14662 17436
rect 14686 17434 14742 17436
rect 14766 17434 14822 17436
rect 14526 17382 14552 17434
rect 14552 17382 14582 17434
rect 14606 17382 14616 17434
rect 14616 17382 14662 17434
rect 14686 17382 14732 17434
rect 14732 17382 14742 17434
rect 14766 17382 14796 17434
rect 14796 17382 14822 17434
rect 14526 17380 14582 17382
rect 14606 17380 14662 17382
rect 14686 17380 14742 17382
rect 14766 17380 14822 17382
rect 14526 16346 14582 16348
rect 14606 16346 14662 16348
rect 14686 16346 14742 16348
rect 14766 16346 14822 16348
rect 14526 16294 14552 16346
rect 14552 16294 14582 16346
rect 14606 16294 14616 16346
rect 14616 16294 14662 16346
rect 14686 16294 14732 16346
rect 14732 16294 14742 16346
rect 14766 16294 14796 16346
rect 14796 16294 14822 16346
rect 14526 16292 14582 16294
rect 14606 16292 14662 16294
rect 14686 16292 14742 16294
rect 14766 16292 14822 16294
rect 14526 15258 14582 15260
rect 14606 15258 14662 15260
rect 14686 15258 14742 15260
rect 14766 15258 14822 15260
rect 14526 15206 14552 15258
rect 14552 15206 14582 15258
rect 14606 15206 14616 15258
rect 14616 15206 14662 15258
rect 14686 15206 14732 15258
rect 14732 15206 14742 15258
rect 14766 15206 14796 15258
rect 14796 15206 14822 15258
rect 14526 15204 14582 15206
rect 14606 15204 14662 15206
rect 14686 15204 14742 15206
rect 14766 15204 14822 15206
rect 16394 15000 16450 15056
rect 14526 14170 14582 14172
rect 14606 14170 14662 14172
rect 14686 14170 14742 14172
rect 14766 14170 14822 14172
rect 14526 14118 14552 14170
rect 14552 14118 14582 14170
rect 14606 14118 14616 14170
rect 14616 14118 14662 14170
rect 14686 14118 14732 14170
rect 14732 14118 14742 14170
rect 14766 14118 14796 14170
rect 14796 14118 14822 14170
rect 14526 14116 14582 14118
rect 14606 14116 14662 14118
rect 14686 14116 14742 14118
rect 14766 14116 14822 14118
rect 14526 13082 14582 13084
rect 14606 13082 14662 13084
rect 14686 13082 14742 13084
rect 14766 13082 14822 13084
rect 14526 13030 14552 13082
rect 14552 13030 14582 13082
rect 14606 13030 14616 13082
rect 14616 13030 14662 13082
rect 14686 13030 14732 13082
rect 14732 13030 14742 13082
rect 14766 13030 14796 13082
rect 14796 13030 14822 13082
rect 14526 13028 14582 13030
rect 14606 13028 14662 13030
rect 14686 13028 14742 13030
rect 14766 13028 14822 13030
rect 14526 11994 14582 11996
rect 14606 11994 14662 11996
rect 14686 11994 14742 11996
rect 14766 11994 14822 11996
rect 14526 11942 14552 11994
rect 14552 11942 14582 11994
rect 14606 11942 14616 11994
rect 14616 11942 14662 11994
rect 14686 11942 14732 11994
rect 14732 11942 14742 11994
rect 14766 11942 14796 11994
rect 14796 11942 14822 11994
rect 14526 11940 14582 11942
rect 14606 11940 14662 11942
rect 14686 11940 14742 11942
rect 14766 11940 14822 11942
rect 15106 12280 15162 12336
rect 9098 7642 9154 7644
rect 9178 7642 9234 7644
rect 9258 7642 9314 7644
rect 9338 7642 9394 7644
rect 9098 7590 9124 7642
rect 9124 7590 9154 7642
rect 9178 7590 9188 7642
rect 9188 7590 9234 7642
rect 9258 7590 9304 7642
rect 9304 7590 9314 7642
rect 9338 7590 9368 7642
rect 9368 7590 9394 7642
rect 9098 7588 9154 7590
rect 9178 7588 9234 7590
rect 9258 7588 9314 7590
rect 9338 7588 9394 7590
rect 9098 6554 9154 6556
rect 9178 6554 9234 6556
rect 9258 6554 9314 6556
rect 9338 6554 9394 6556
rect 9098 6502 9124 6554
rect 9124 6502 9154 6554
rect 9178 6502 9188 6554
rect 9188 6502 9234 6554
rect 9258 6502 9304 6554
rect 9304 6502 9314 6554
rect 9338 6502 9368 6554
rect 9368 6502 9394 6554
rect 9098 6500 9154 6502
rect 9178 6500 9234 6502
rect 9258 6500 9314 6502
rect 9338 6500 9394 6502
rect 9098 5466 9154 5468
rect 9178 5466 9234 5468
rect 9258 5466 9314 5468
rect 9338 5466 9394 5468
rect 9098 5414 9124 5466
rect 9124 5414 9154 5466
rect 9178 5414 9188 5466
rect 9188 5414 9234 5466
rect 9258 5414 9304 5466
rect 9304 5414 9314 5466
rect 9338 5414 9368 5466
rect 9368 5414 9394 5466
rect 9098 5412 9154 5414
rect 9178 5412 9234 5414
rect 9258 5412 9314 5414
rect 9338 5412 9394 5414
rect 9098 4378 9154 4380
rect 9178 4378 9234 4380
rect 9258 4378 9314 4380
rect 9338 4378 9394 4380
rect 9098 4326 9124 4378
rect 9124 4326 9154 4378
rect 9178 4326 9188 4378
rect 9188 4326 9234 4378
rect 9258 4326 9304 4378
rect 9304 4326 9314 4378
rect 9338 4326 9368 4378
rect 9368 4326 9394 4378
rect 9098 4324 9154 4326
rect 9178 4324 9234 4326
rect 9258 4324 9314 4326
rect 9338 4324 9394 4326
rect 11812 9274 11868 9276
rect 11892 9274 11948 9276
rect 11972 9274 12028 9276
rect 12052 9274 12108 9276
rect 11812 9222 11838 9274
rect 11838 9222 11868 9274
rect 11892 9222 11902 9274
rect 11902 9222 11948 9274
rect 11972 9222 12018 9274
rect 12018 9222 12028 9274
rect 12052 9222 12082 9274
rect 12082 9222 12108 9274
rect 11812 9220 11868 9222
rect 11892 9220 11948 9222
rect 11972 9220 12028 9222
rect 12052 9220 12108 9222
rect 11812 8186 11868 8188
rect 11892 8186 11948 8188
rect 11972 8186 12028 8188
rect 12052 8186 12108 8188
rect 11812 8134 11838 8186
rect 11838 8134 11868 8186
rect 11892 8134 11902 8186
rect 11902 8134 11948 8186
rect 11972 8134 12018 8186
rect 12018 8134 12028 8186
rect 12052 8134 12082 8186
rect 12082 8134 12108 8186
rect 11812 8132 11868 8134
rect 11892 8132 11948 8134
rect 11972 8132 12028 8134
rect 12052 8132 12108 8134
rect 11812 7098 11868 7100
rect 11892 7098 11948 7100
rect 11972 7098 12028 7100
rect 12052 7098 12108 7100
rect 11812 7046 11838 7098
rect 11838 7046 11868 7098
rect 11892 7046 11902 7098
rect 11902 7046 11948 7098
rect 11972 7046 12018 7098
rect 12018 7046 12028 7098
rect 12052 7046 12082 7098
rect 12082 7046 12108 7098
rect 11812 7044 11868 7046
rect 11892 7044 11948 7046
rect 11972 7044 12028 7046
rect 12052 7044 12108 7046
rect 14526 10906 14582 10908
rect 14606 10906 14662 10908
rect 14686 10906 14742 10908
rect 14766 10906 14822 10908
rect 14526 10854 14552 10906
rect 14552 10854 14582 10906
rect 14606 10854 14616 10906
rect 14616 10854 14662 10906
rect 14686 10854 14732 10906
rect 14732 10854 14742 10906
rect 14766 10854 14796 10906
rect 14796 10854 14822 10906
rect 14526 10852 14582 10854
rect 14606 10852 14662 10854
rect 14686 10852 14742 10854
rect 14766 10852 14822 10854
rect 14526 9818 14582 9820
rect 14606 9818 14662 9820
rect 14686 9818 14742 9820
rect 14766 9818 14822 9820
rect 14526 9766 14552 9818
rect 14552 9766 14582 9818
rect 14606 9766 14616 9818
rect 14616 9766 14662 9818
rect 14686 9766 14732 9818
rect 14732 9766 14742 9818
rect 14766 9766 14796 9818
rect 14796 9766 14822 9818
rect 14526 9764 14582 9766
rect 14606 9764 14662 9766
rect 14686 9764 14742 9766
rect 14766 9764 14822 9766
rect 11812 6010 11868 6012
rect 11892 6010 11948 6012
rect 11972 6010 12028 6012
rect 12052 6010 12108 6012
rect 11812 5958 11838 6010
rect 11838 5958 11868 6010
rect 11892 5958 11902 6010
rect 11902 5958 11948 6010
rect 11972 5958 12018 6010
rect 12018 5958 12028 6010
rect 12052 5958 12082 6010
rect 12082 5958 12108 6010
rect 11812 5956 11868 5958
rect 11892 5956 11948 5958
rect 11972 5956 12028 5958
rect 12052 5956 12108 5958
rect 6384 2746 6440 2748
rect 6464 2746 6520 2748
rect 6544 2746 6600 2748
rect 6624 2746 6680 2748
rect 6384 2694 6410 2746
rect 6410 2694 6440 2746
rect 6464 2694 6474 2746
rect 6474 2694 6520 2746
rect 6544 2694 6590 2746
rect 6590 2694 6600 2746
rect 6624 2694 6654 2746
rect 6654 2694 6680 2746
rect 6384 2692 6440 2694
rect 6464 2692 6520 2694
rect 6544 2692 6600 2694
rect 6624 2692 6680 2694
rect 9098 3290 9154 3292
rect 9178 3290 9234 3292
rect 9258 3290 9314 3292
rect 9338 3290 9394 3292
rect 9098 3238 9124 3290
rect 9124 3238 9154 3290
rect 9178 3238 9188 3290
rect 9188 3238 9234 3290
rect 9258 3238 9304 3290
rect 9304 3238 9314 3290
rect 9338 3238 9368 3290
rect 9368 3238 9394 3290
rect 9098 3236 9154 3238
rect 9178 3236 9234 3238
rect 9258 3236 9314 3238
rect 9338 3236 9394 3238
rect 9098 2202 9154 2204
rect 9178 2202 9234 2204
rect 9258 2202 9314 2204
rect 9338 2202 9394 2204
rect 9098 2150 9124 2202
rect 9124 2150 9154 2202
rect 9178 2150 9188 2202
rect 9188 2150 9234 2202
rect 9258 2150 9304 2202
rect 9304 2150 9314 2202
rect 9338 2150 9368 2202
rect 9368 2150 9394 2202
rect 9098 2148 9154 2150
rect 9178 2148 9234 2150
rect 9258 2148 9314 2150
rect 9338 2148 9394 2150
rect 11812 4922 11868 4924
rect 11892 4922 11948 4924
rect 11972 4922 12028 4924
rect 12052 4922 12108 4924
rect 11812 4870 11838 4922
rect 11838 4870 11868 4922
rect 11892 4870 11902 4922
rect 11902 4870 11948 4922
rect 11972 4870 12018 4922
rect 12018 4870 12028 4922
rect 12052 4870 12082 4922
rect 12082 4870 12108 4922
rect 11812 4868 11868 4870
rect 11892 4868 11948 4870
rect 11972 4868 12028 4870
rect 12052 4868 12108 4870
rect 11812 3834 11868 3836
rect 11892 3834 11948 3836
rect 11972 3834 12028 3836
rect 12052 3834 12108 3836
rect 11812 3782 11838 3834
rect 11838 3782 11868 3834
rect 11892 3782 11902 3834
rect 11902 3782 11948 3834
rect 11972 3782 12018 3834
rect 12018 3782 12028 3834
rect 12052 3782 12082 3834
rect 12082 3782 12108 3834
rect 11812 3780 11868 3782
rect 11892 3780 11948 3782
rect 11972 3780 12028 3782
rect 12052 3780 12108 3782
rect 11812 2746 11868 2748
rect 11892 2746 11948 2748
rect 11972 2746 12028 2748
rect 12052 2746 12108 2748
rect 11812 2694 11838 2746
rect 11838 2694 11868 2746
rect 11892 2694 11902 2746
rect 11902 2694 11948 2746
rect 11972 2694 12018 2746
rect 12018 2694 12028 2746
rect 12052 2694 12082 2746
rect 12082 2694 12108 2746
rect 11812 2692 11868 2694
rect 11892 2692 11948 2694
rect 11972 2692 12028 2694
rect 12052 2692 12108 2694
rect 14526 8730 14582 8732
rect 14606 8730 14662 8732
rect 14686 8730 14742 8732
rect 14766 8730 14822 8732
rect 14526 8678 14552 8730
rect 14552 8678 14582 8730
rect 14606 8678 14616 8730
rect 14616 8678 14662 8730
rect 14686 8678 14732 8730
rect 14732 8678 14742 8730
rect 14766 8678 14796 8730
rect 14796 8678 14822 8730
rect 14526 8676 14582 8678
rect 14606 8676 14662 8678
rect 14686 8676 14742 8678
rect 14766 8676 14822 8678
rect 14526 7642 14582 7644
rect 14606 7642 14662 7644
rect 14686 7642 14742 7644
rect 14766 7642 14822 7644
rect 14526 7590 14552 7642
rect 14552 7590 14582 7642
rect 14606 7590 14616 7642
rect 14616 7590 14662 7642
rect 14686 7590 14732 7642
rect 14732 7590 14742 7642
rect 14766 7590 14796 7642
rect 14796 7590 14822 7642
rect 14526 7588 14582 7590
rect 14606 7588 14662 7590
rect 14686 7588 14742 7590
rect 14766 7588 14822 7590
rect 14526 6554 14582 6556
rect 14606 6554 14662 6556
rect 14686 6554 14742 6556
rect 14766 6554 14822 6556
rect 14526 6502 14552 6554
rect 14552 6502 14582 6554
rect 14606 6502 14616 6554
rect 14616 6502 14662 6554
rect 14686 6502 14732 6554
rect 14732 6502 14742 6554
rect 14766 6502 14796 6554
rect 14796 6502 14822 6554
rect 14526 6500 14582 6502
rect 14606 6500 14662 6502
rect 14686 6500 14742 6502
rect 14766 6500 14822 6502
rect 16394 9560 16450 9616
rect 16670 7520 16726 7576
rect 14526 5466 14582 5468
rect 14606 5466 14662 5468
rect 14686 5466 14742 5468
rect 14766 5466 14822 5468
rect 14526 5414 14552 5466
rect 14552 5414 14582 5466
rect 14606 5414 14616 5466
rect 14616 5414 14662 5466
rect 14686 5414 14732 5466
rect 14732 5414 14742 5466
rect 14766 5414 14796 5466
rect 14796 5414 14822 5466
rect 14526 5412 14582 5414
rect 14606 5412 14662 5414
rect 14686 5412 14742 5414
rect 14766 5412 14822 5414
rect 14526 4378 14582 4380
rect 14606 4378 14662 4380
rect 14686 4378 14742 4380
rect 14766 4378 14822 4380
rect 14526 4326 14552 4378
rect 14552 4326 14582 4378
rect 14606 4326 14616 4378
rect 14616 4326 14662 4378
rect 14686 4326 14732 4378
rect 14732 4326 14742 4378
rect 14766 4326 14796 4378
rect 14796 4326 14822 4378
rect 14526 4324 14582 4326
rect 14606 4324 14662 4326
rect 14686 4324 14742 4326
rect 14766 4324 14822 4326
rect 14526 3290 14582 3292
rect 14606 3290 14662 3292
rect 14686 3290 14742 3292
rect 14766 3290 14822 3292
rect 14526 3238 14552 3290
rect 14552 3238 14582 3290
rect 14606 3238 14616 3290
rect 14616 3238 14662 3290
rect 14686 3238 14732 3290
rect 14732 3238 14742 3290
rect 14766 3238 14796 3290
rect 14796 3238 14822 3290
rect 14526 3236 14582 3238
rect 14606 3236 14662 3238
rect 14686 3236 14742 3238
rect 14766 3236 14822 3238
rect 14526 2202 14582 2204
rect 14606 2202 14662 2204
rect 14686 2202 14742 2204
rect 14766 2202 14822 2204
rect 14526 2150 14552 2202
rect 14552 2150 14582 2202
rect 14606 2150 14616 2202
rect 14616 2150 14662 2202
rect 14686 2150 14732 2202
rect 14732 2150 14742 2202
rect 14766 2150 14796 2202
rect 14796 2150 14822 2202
rect 14526 2148 14582 2150
rect 14606 2148 14662 2150
rect 14686 2148 14742 2150
rect 14766 2148 14822 2150
rect 16394 4800 16450 4856
rect 15750 2080 15806 2136
<< metal3 >>
rect 3658 18528 3978 18529
rect 0 18458 800 18488
rect 3658 18464 3666 18528
rect 3730 18464 3746 18528
rect 3810 18464 3826 18528
rect 3890 18464 3906 18528
rect 3970 18464 3978 18528
rect 3658 18463 3978 18464
rect 9086 18528 9406 18529
rect 9086 18464 9094 18528
rect 9158 18464 9174 18528
rect 9238 18464 9254 18528
rect 9318 18464 9334 18528
rect 9398 18464 9406 18528
rect 9086 18463 9406 18464
rect 14514 18528 14834 18529
rect 14514 18464 14522 18528
rect 14586 18464 14602 18528
rect 14666 18464 14682 18528
rect 14746 18464 14762 18528
rect 14826 18464 14834 18528
rect 14514 18463 14834 18464
rect 1761 18458 1827 18461
rect 0 18456 1827 18458
rect 0 18400 1766 18456
rect 1822 18400 1827 18456
rect 0 18398 1827 18400
rect 0 18368 800 18398
rect 1761 18395 1827 18398
rect 6372 17984 6692 17985
rect 6372 17920 6380 17984
rect 6444 17920 6460 17984
rect 6524 17920 6540 17984
rect 6604 17920 6620 17984
rect 6684 17920 6692 17984
rect 6372 17919 6692 17920
rect 11800 17984 12120 17985
rect 11800 17920 11808 17984
rect 11872 17920 11888 17984
rect 11952 17920 11968 17984
rect 12032 17920 12048 17984
rect 12112 17920 12120 17984
rect 11800 17919 12120 17920
rect 13813 17778 13879 17781
rect 17748 17778 18548 17808
rect 13813 17776 18548 17778
rect 13813 17720 13818 17776
rect 13874 17720 18548 17776
rect 13813 17718 18548 17720
rect 13813 17715 13879 17718
rect 17748 17688 18548 17718
rect 3658 17440 3978 17441
rect 3658 17376 3666 17440
rect 3730 17376 3746 17440
rect 3810 17376 3826 17440
rect 3890 17376 3906 17440
rect 3970 17376 3978 17440
rect 3658 17375 3978 17376
rect 9086 17440 9406 17441
rect 9086 17376 9094 17440
rect 9158 17376 9174 17440
rect 9238 17376 9254 17440
rect 9318 17376 9334 17440
rect 9398 17376 9406 17440
rect 9086 17375 9406 17376
rect 14514 17440 14834 17441
rect 14514 17376 14522 17440
rect 14586 17376 14602 17440
rect 14666 17376 14682 17440
rect 14746 17376 14762 17440
rect 14826 17376 14834 17440
rect 14514 17375 14834 17376
rect 6372 16896 6692 16897
rect 6372 16832 6380 16896
rect 6444 16832 6460 16896
rect 6524 16832 6540 16896
rect 6604 16832 6620 16896
rect 6684 16832 6692 16896
rect 6372 16831 6692 16832
rect 11800 16896 12120 16897
rect 11800 16832 11808 16896
rect 11872 16832 11888 16896
rect 11952 16832 11968 16896
rect 12032 16832 12048 16896
rect 12112 16832 12120 16896
rect 11800 16831 12120 16832
rect 3658 16352 3978 16353
rect 3658 16288 3666 16352
rect 3730 16288 3746 16352
rect 3810 16288 3826 16352
rect 3890 16288 3906 16352
rect 3970 16288 3978 16352
rect 3658 16287 3978 16288
rect 9086 16352 9406 16353
rect 9086 16288 9094 16352
rect 9158 16288 9174 16352
rect 9238 16288 9254 16352
rect 9318 16288 9334 16352
rect 9398 16288 9406 16352
rect 9086 16287 9406 16288
rect 14514 16352 14834 16353
rect 14514 16288 14522 16352
rect 14586 16288 14602 16352
rect 14666 16288 14682 16352
rect 14746 16288 14762 16352
rect 14826 16288 14834 16352
rect 14514 16287 14834 16288
rect 6372 15808 6692 15809
rect 0 15738 800 15768
rect 6372 15744 6380 15808
rect 6444 15744 6460 15808
rect 6524 15744 6540 15808
rect 6604 15744 6620 15808
rect 6684 15744 6692 15808
rect 6372 15743 6692 15744
rect 11800 15808 12120 15809
rect 11800 15744 11808 15808
rect 11872 15744 11888 15808
rect 11952 15744 11968 15808
rect 12032 15744 12048 15808
rect 12112 15744 12120 15808
rect 11800 15743 12120 15744
rect 1945 15738 2011 15741
rect 0 15736 2011 15738
rect 0 15680 1950 15736
rect 2006 15680 2011 15736
rect 0 15678 2011 15680
rect 0 15648 800 15678
rect 1945 15675 2011 15678
rect 3658 15264 3978 15265
rect 3658 15200 3666 15264
rect 3730 15200 3746 15264
rect 3810 15200 3826 15264
rect 3890 15200 3906 15264
rect 3970 15200 3978 15264
rect 3658 15199 3978 15200
rect 9086 15264 9406 15265
rect 9086 15200 9094 15264
rect 9158 15200 9174 15264
rect 9238 15200 9254 15264
rect 9318 15200 9334 15264
rect 9398 15200 9406 15264
rect 9086 15199 9406 15200
rect 14514 15264 14834 15265
rect 14514 15200 14522 15264
rect 14586 15200 14602 15264
rect 14666 15200 14682 15264
rect 14746 15200 14762 15264
rect 14826 15200 14834 15264
rect 14514 15199 14834 15200
rect 16389 15058 16455 15061
rect 17748 15058 18548 15088
rect 16389 15056 18548 15058
rect 16389 15000 16394 15056
rect 16450 15000 18548 15056
rect 16389 14998 18548 15000
rect 16389 14995 16455 14998
rect 17748 14968 18548 14998
rect 6372 14720 6692 14721
rect 6372 14656 6380 14720
rect 6444 14656 6460 14720
rect 6524 14656 6540 14720
rect 6604 14656 6620 14720
rect 6684 14656 6692 14720
rect 6372 14655 6692 14656
rect 11800 14720 12120 14721
rect 11800 14656 11808 14720
rect 11872 14656 11888 14720
rect 11952 14656 11968 14720
rect 12032 14656 12048 14720
rect 12112 14656 12120 14720
rect 11800 14655 12120 14656
rect 3658 14176 3978 14177
rect 3658 14112 3666 14176
rect 3730 14112 3746 14176
rect 3810 14112 3826 14176
rect 3890 14112 3906 14176
rect 3970 14112 3978 14176
rect 3658 14111 3978 14112
rect 9086 14176 9406 14177
rect 9086 14112 9094 14176
rect 9158 14112 9174 14176
rect 9238 14112 9254 14176
rect 9318 14112 9334 14176
rect 9398 14112 9406 14176
rect 9086 14111 9406 14112
rect 14514 14176 14834 14177
rect 14514 14112 14522 14176
rect 14586 14112 14602 14176
rect 14666 14112 14682 14176
rect 14746 14112 14762 14176
rect 14826 14112 14834 14176
rect 14514 14111 14834 14112
rect 6372 13632 6692 13633
rect 6372 13568 6380 13632
rect 6444 13568 6460 13632
rect 6524 13568 6540 13632
rect 6604 13568 6620 13632
rect 6684 13568 6692 13632
rect 6372 13567 6692 13568
rect 11800 13632 12120 13633
rect 11800 13568 11808 13632
rect 11872 13568 11888 13632
rect 11952 13568 11968 13632
rect 12032 13568 12048 13632
rect 12112 13568 12120 13632
rect 11800 13567 12120 13568
rect 3658 13088 3978 13089
rect 0 13018 800 13048
rect 3658 13024 3666 13088
rect 3730 13024 3746 13088
rect 3810 13024 3826 13088
rect 3890 13024 3906 13088
rect 3970 13024 3978 13088
rect 3658 13023 3978 13024
rect 9086 13088 9406 13089
rect 9086 13024 9094 13088
rect 9158 13024 9174 13088
rect 9238 13024 9254 13088
rect 9318 13024 9334 13088
rect 9398 13024 9406 13088
rect 9086 13023 9406 13024
rect 14514 13088 14834 13089
rect 14514 13024 14522 13088
rect 14586 13024 14602 13088
rect 14666 13024 14682 13088
rect 14746 13024 14762 13088
rect 14826 13024 14834 13088
rect 14514 13023 14834 13024
rect 2773 13018 2839 13021
rect 0 13016 2839 13018
rect 0 12960 2778 13016
rect 2834 12960 2839 13016
rect 0 12958 2839 12960
rect 0 12928 800 12958
rect 2773 12955 2839 12958
rect 6372 12544 6692 12545
rect 6372 12480 6380 12544
rect 6444 12480 6460 12544
rect 6524 12480 6540 12544
rect 6604 12480 6620 12544
rect 6684 12480 6692 12544
rect 6372 12479 6692 12480
rect 11800 12544 12120 12545
rect 11800 12480 11808 12544
rect 11872 12480 11888 12544
rect 11952 12480 11968 12544
rect 12032 12480 12048 12544
rect 12112 12480 12120 12544
rect 11800 12479 12120 12480
rect 15101 12338 15167 12341
rect 17748 12338 18548 12368
rect 15101 12336 18548 12338
rect 15101 12280 15106 12336
rect 15162 12280 18548 12336
rect 15101 12278 18548 12280
rect 15101 12275 15167 12278
rect 17748 12248 18548 12278
rect 3658 12000 3978 12001
rect 3658 11936 3666 12000
rect 3730 11936 3746 12000
rect 3810 11936 3826 12000
rect 3890 11936 3906 12000
rect 3970 11936 3978 12000
rect 3658 11935 3978 11936
rect 9086 12000 9406 12001
rect 9086 11936 9094 12000
rect 9158 11936 9174 12000
rect 9238 11936 9254 12000
rect 9318 11936 9334 12000
rect 9398 11936 9406 12000
rect 9086 11935 9406 11936
rect 14514 12000 14834 12001
rect 14514 11936 14522 12000
rect 14586 11936 14602 12000
rect 14666 11936 14682 12000
rect 14746 11936 14762 12000
rect 14826 11936 14834 12000
rect 14514 11935 14834 11936
rect 6372 11456 6692 11457
rect 6372 11392 6380 11456
rect 6444 11392 6460 11456
rect 6524 11392 6540 11456
rect 6604 11392 6620 11456
rect 6684 11392 6692 11456
rect 6372 11391 6692 11392
rect 11800 11456 12120 11457
rect 11800 11392 11808 11456
rect 11872 11392 11888 11456
rect 11952 11392 11968 11456
rect 12032 11392 12048 11456
rect 12112 11392 12120 11456
rect 11800 11391 12120 11392
rect 0 10978 800 11008
rect 1761 10978 1827 10981
rect 0 10976 1827 10978
rect 0 10920 1766 10976
rect 1822 10920 1827 10976
rect 0 10918 1827 10920
rect 0 10888 800 10918
rect 1761 10915 1827 10918
rect 3658 10912 3978 10913
rect 3658 10848 3666 10912
rect 3730 10848 3746 10912
rect 3810 10848 3826 10912
rect 3890 10848 3906 10912
rect 3970 10848 3978 10912
rect 3658 10847 3978 10848
rect 9086 10912 9406 10913
rect 9086 10848 9094 10912
rect 9158 10848 9174 10912
rect 9238 10848 9254 10912
rect 9318 10848 9334 10912
rect 9398 10848 9406 10912
rect 9086 10847 9406 10848
rect 14514 10912 14834 10913
rect 14514 10848 14522 10912
rect 14586 10848 14602 10912
rect 14666 10848 14682 10912
rect 14746 10848 14762 10912
rect 14826 10848 14834 10912
rect 14514 10847 14834 10848
rect 6372 10368 6692 10369
rect 6372 10304 6380 10368
rect 6444 10304 6460 10368
rect 6524 10304 6540 10368
rect 6604 10304 6620 10368
rect 6684 10304 6692 10368
rect 6372 10303 6692 10304
rect 11800 10368 12120 10369
rect 11800 10304 11808 10368
rect 11872 10304 11888 10368
rect 11952 10304 11968 10368
rect 12032 10304 12048 10368
rect 12112 10304 12120 10368
rect 11800 10303 12120 10304
rect 3658 9824 3978 9825
rect 3658 9760 3666 9824
rect 3730 9760 3746 9824
rect 3810 9760 3826 9824
rect 3890 9760 3906 9824
rect 3970 9760 3978 9824
rect 3658 9759 3978 9760
rect 9086 9824 9406 9825
rect 9086 9760 9094 9824
rect 9158 9760 9174 9824
rect 9238 9760 9254 9824
rect 9318 9760 9334 9824
rect 9398 9760 9406 9824
rect 9086 9759 9406 9760
rect 14514 9824 14834 9825
rect 14514 9760 14522 9824
rect 14586 9760 14602 9824
rect 14666 9760 14682 9824
rect 14746 9760 14762 9824
rect 14826 9760 14834 9824
rect 14514 9759 14834 9760
rect 4705 9618 4771 9621
rect 8569 9618 8635 9621
rect 4705 9616 8635 9618
rect 4705 9560 4710 9616
rect 4766 9560 8574 9616
rect 8630 9560 8635 9616
rect 4705 9558 8635 9560
rect 4705 9555 4771 9558
rect 8569 9555 8635 9558
rect 16389 9618 16455 9621
rect 17748 9618 18548 9648
rect 16389 9616 18548 9618
rect 16389 9560 16394 9616
rect 16450 9560 18548 9616
rect 16389 9558 18548 9560
rect 16389 9555 16455 9558
rect 17748 9528 18548 9558
rect 6372 9280 6692 9281
rect 6372 9216 6380 9280
rect 6444 9216 6460 9280
rect 6524 9216 6540 9280
rect 6604 9216 6620 9280
rect 6684 9216 6692 9280
rect 6372 9215 6692 9216
rect 11800 9280 12120 9281
rect 11800 9216 11808 9280
rect 11872 9216 11888 9280
rect 11952 9216 11968 9280
rect 12032 9216 12048 9280
rect 12112 9216 12120 9280
rect 11800 9215 12120 9216
rect 3658 8736 3978 8737
rect 3658 8672 3666 8736
rect 3730 8672 3746 8736
rect 3810 8672 3826 8736
rect 3890 8672 3906 8736
rect 3970 8672 3978 8736
rect 3658 8671 3978 8672
rect 9086 8736 9406 8737
rect 9086 8672 9094 8736
rect 9158 8672 9174 8736
rect 9238 8672 9254 8736
rect 9318 8672 9334 8736
rect 9398 8672 9406 8736
rect 9086 8671 9406 8672
rect 14514 8736 14834 8737
rect 14514 8672 14522 8736
rect 14586 8672 14602 8736
rect 14666 8672 14682 8736
rect 14746 8672 14762 8736
rect 14826 8672 14834 8736
rect 14514 8671 14834 8672
rect 0 8258 800 8288
rect 1945 8258 2011 8261
rect 0 8256 2011 8258
rect 0 8200 1950 8256
rect 2006 8200 2011 8256
rect 0 8198 2011 8200
rect 0 8168 800 8198
rect 1945 8195 2011 8198
rect 6372 8192 6692 8193
rect 6372 8128 6380 8192
rect 6444 8128 6460 8192
rect 6524 8128 6540 8192
rect 6604 8128 6620 8192
rect 6684 8128 6692 8192
rect 6372 8127 6692 8128
rect 11800 8192 12120 8193
rect 11800 8128 11808 8192
rect 11872 8128 11888 8192
rect 11952 8128 11968 8192
rect 12032 8128 12048 8192
rect 12112 8128 12120 8192
rect 11800 8127 12120 8128
rect 3658 7648 3978 7649
rect 3658 7584 3666 7648
rect 3730 7584 3746 7648
rect 3810 7584 3826 7648
rect 3890 7584 3906 7648
rect 3970 7584 3978 7648
rect 3658 7583 3978 7584
rect 9086 7648 9406 7649
rect 9086 7584 9094 7648
rect 9158 7584 9174 7648
rect 9238 7584 9254 7648
rect 9318 7584 9334 7648
rect 9398 7584 9406 7648
rect 9086 7583 9406 7584
rect 14514 7648 14834 7649
rect 14514 7584 14522 7648
rect 14586 7584 14602 7648
rect 14666 7584 14682 7648
rect 14746 7584 14762 7648
rect 14826 7584 14834 7648
rect 14514 7583 14834 7584
rect 16665 7578 16731 7581
rect 17748 7578 18548 7608
rect 16665 7576 18548 7578
rect 16665 7520 16670 7576
rect 16726 7520 18548 7576
rect 16665 7518 18548 7520
rect 16665 7515 16731 7518
rect 17748 7488 18548 7518
rect 6372 7104 6692 7105
rect 6372 7040 6380 7104
rect 6444 7040 6460 7104
rect 6524 7040 6540 7104
rect 6604 7040 6620 7104
rect 6684 7040 6692 7104
rect 6372 7039 6692 7040
rect 11800 7104 12120 7105
rect 11800 7040 11808 7104
rect 11872 7040 11888 7104
rect 11952 7040 11968 7104
rect 12032 7040 12048 7104
rect 12112 7040 12120 7104
rect 11800 7039 12120 7040
rect 3658 6560 3978 6561
rect 3658 6496 3666 6560
rect 3730 6496 3746 6560
rect 3810 6496 3826 6560
rect 3890 6496 3906 6560
rect 3970 6496 3978 6560
rect 3658 6495 3978 6496
rect 9086 6560 9406 6561
rect 9086 6496 9094 6560
rect 9158 6496 9174 6560
rect 9238 6496 9254 6560
rect 9318 6496 9334 6560
rect 9398 6496 9406 6560
rect 9086 6495 9406 6496
rect 14514 6560 14834 6561
rect 14514 6496 14522 6560
rect 14586 6496 14602 6560
rect 14666 6496 14682 6560
rect 14746 6496 14762 6560
rect 14826 6496 14834 6560
rect 14514 6495 14834 6496
rect 6372 6016 6692 6017
rect 6372 5952 6380 6016
rect 6444 5952 6460 6016
rect 6524 5952 6540 6016
rect 6604 5952 6620 6016
rect 6684 5952 6692 6016
rect 6372 5951 6692 5952
rect 11800 6016 12120 6017
rect 11800 5952 11808 6016
rect 11872 5952 11888 6016
rect 11952 5952 11968 6016
rect 12032 5952 12048 6016
rect 12112 5952 12120 6016
rect 11800 5951 12120 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 3658 5472 3978 5473
rect 3658 5408 3666 5472
rect 3730 5408 3746 5472
rect 3810 5408 3826 5472
rect 3890 5408 3906 5472
rect 3970 5408 3978 5472
rect 3658 5407 3978 5408
rect 9086 5472 9406 5473
rect 9086 5408 9094 5472
rect 9158 5408 9174 5472
rect 9238 5408 9254 5472
rect 9318 5408 9334 5472
rect 9398 5408 9406 5472
rect 9086 5407 9406 5408
rect 14514 5472 14834 5473
rect 14514 5408 14522 5472
rect 14586 5408 14602 5472
rect 14666 5408 14682 5472
rect 14746 5408 14762 5472
rect 14826 5408 14834 5472
rect 14514 5407 14834 5408
rect 6372 4928 6692 4929
rect 6372 4864 6380 4928
rect 6444 4864 6460 4928
rect 6524 4864 6540 4928
rect 6604 4864 6620 4928
rect 6684 4864 6692 4928
rect 6372 4863 6692 4864
rect 11800 4928 12120 4929
rect 11800 4864 11808 4928
rect 11872 4864 11888 4928
rect 11952 4864 11968 4928
rect 12032 4864 12048 4928
rect 12112 4864 12120 4928
rect 11800 4863 12120 4864
rect 16389 4858 16455 4861
rect 17748 4858 18548 4888
rect 16389 4856 18548 4858
rect 16389 4800 16394 4856
rect 16450 4800 18548 4856
rect 16389 4798 18548 4800
rect 16389 4795 16455 4798
rect 17748 4768 18548 4798
rect 3658 4384 3978 4385
rect 3658 4320 3666 4384
rect 3730 4320 3746 4384
rect 3810 4320 3826 4384
rect 3890 4320 3906 4384
rect 3970 4320 3978 4384
rect 3658 4319 3978 4320
rect 9086 4384 9406 4385
rect 9086 4320 9094 4384
rect 9158 4320 9174 4384
rect 9238 4320 9254 4384
rect 9318 4320 9334 4384
rect 9398 4320 9406 4384
rect 9086 4319 9406 4320
rect 14514 4384 14834 4385
rect 14514 4320 14522 4384
rect 14586 4320 14602 4384
rect 14666 4320 14682 4384
rect 14746 4320 14762 4384
rect 14826 4320 14834 4384
rect 14514 4319 14834 4320
rect 6372 3840 6692 3841
rect 6372 3776 6380 3840
rect 6444 3776 6460 3840
rect 6524 3776 6540 3840
rect 6604 3776 6620 3840
rect 6684 3776 6692 3840
rect 6372 3775 6692 3776
rect 11800 3840 12120 3841
rect 11800 3776 11808 3840
rect 11872 3776 11888 3840
rect 11952 3776 11968 3840
rect 12032 3776 12048 3840
rect 12112 3776 12120 3840
rect 11800 3775 12120 3776
rect 3658 3296 3978 3297
rect 3658 3232 3666 3296
rect 3730 3232 3746 3296
rect 3810 3232 3826 3296
rect 3890 3232 3906 3296
rect 3970 3232 3978 3296
rect 3658 3231 3978 3232
rect 9086 3296 9406 3297
rect 9086 3232 9094 3296
rect 9158 3232 9174 3296
rect 9238 3232 9254 3296
rect 9318 3232 9334 3296
rect 9398 3232 9406 3296
rect 9086 3231 9406 3232
rect 14514 3296 14834 3297
rect 14514 3232 14522 3296
rect 14586 3232 14602 3296
rect 14666 3232 14682 3296
rect 14746 3232 14762 3296
rect 14826 3232 14834 3296
rect 14514 3231 14834 3232
rect 0 2818 800 2848
rect 3969 2818 4035 2821
rect 0 2816 4035 2818
rect 0 2760 3974 2816
rect 4030 2760 4035 2816
rect 0 2758 4035 2760
rect 0 2728 800 2758
rect 3969 2755 4035 2758
rect 6372 2752 6692 2753
rect 6372 2688 6380 2752
rect 6444 2688 6460 2752
rect 6524 2688 6540 2752
rect 6604 2688 6620 2752
rect 6684 2688 6692 2752
rect 6372 2687 6692 2688
rect 11800 2752 12120 2753
rect 11800 2688 11808 2752
rect 11872 2688 11888 2752
rect 11952 2688 11968 2752
rect 12032 2688 12048 2752
rect 12112 2688 12120 2752
rect 11800 2687 12120 2688
rect 3658 2208 3978 2209
rect 3658 2144 3666 2208
rect 3730 2144 3746 2208
rect 3810 2144 3826 2208
rect 3890 2144 3906 2208
rect 3970 2144 3978 2208
rect 3658 2143 3978 2144
rect 9086 2208 9406 2209
rect 9086 2144 9094 2208
rect 9158 2144 9174 2208
rect 9238 2144 9254 2208
rect 9318 2144 9334 2208
rect 9398 2144 9406 2208
rect 9086 2143 9406 2144
rect 14514 2208 14834 2209
rect 14514 2144 14522 2208
rect 14586 2144 14602 2208
rect 14666 2144 14682 2208
rect 14746 2144 14762 2208
rect 14826 2144 14834 2208
rect 14514 2143 14834 2144
rect 15745 2138 15811 2141
rect 17748 2138 18548 2168
rect 15745 2136 18548 2138
rect 15745 2080 15750 2136
rect 15806 2080 18548 2136
rect 15745 2078 18548 2080
rect 15745 2075 15811 2078
rect 17748 2048 18548 2078
<< via3 >>
rect 3666 18524 3730 18528
rect 3666 18468 3670 18524
rect 3670 18468 3726 18524
rect 3726 18468 3730 18524
rect 3666 18464 3730 18468
rect 3746 18524 3810 18528
rect 3746 18468 3750 18524
rect 3750 18468 3806 18524
rect 3806 18468 3810 18524
rect 3746 18464 3810 18468
rect 3826 18524 3890 18528
rect 3826 18468 3830 18524
rect 3830 18468 3886 18524
rect 3886 18468 3890 18524
rect 3826 18464 3890 18468
rect 3906 18524 3970 18528
rect 3906 18468 3910 18524
rect 3910 18468 3966 18524
rect 3966 18468 3970 18524
rect 3906 18464 3970 18468
rect 9094 18524 9158 18528
rect 9094 18468 9098 18524
rect 9098 18468 9154 18524
rect 9154 18468 9158 18524
rect 9094 18464 9158 18468
rect 9174 18524 9238 18528
rect 9174 18468 9178 18524
rect 9178 18468 9234 18524
rect 9234 18468 9238 18524
rect 9174 18464 9238 18468
rect 9254 18524 9318 18528
rect 9254 18468 9258 18524
rect 9258 18468 9314 18524
rect 9314 18468 9318 18524
rect 9254 18464 9318 18468
rect 9334 18524 9398 18528
rect 9334 18468 9338 18524
rect 9338 18468 9394 18524
rect 9394 18468 9398 18524
rect 9334 18464 9398 18468
rect 14522 18524 14586 18528
rect 14522 18468 14526 18524
rect 14526 18468 14582 18524
rect 14582 18468 14586 18524
rect 14522 18464 14586 18468
rect 14602 18524 14666 18528
rect 14602 18468 14606 18524
rect 14606 18468 14662 18524
rect 14662 18468 14666 18524
rect 14602 18464 14666 18468
rect 14682 18524 14746 18528
rect 14682 18468 14686 18524
rect 14686 18468 14742 18524
rect 14742 18468 14746 18524
rect 14682 18464 14746 18468
rect 14762 18524 14826 18528
rect 14762 18468 14766 18524
rect 14766 18468 14822 18524
rect 14822 18468 14826 18524
rect 14762 18464 14826 18468
rect 6380 17980 6444 17984
rect 6380 17924 6384 17980
rect 6384 17924 6440 17980
rect 6440 17924 6444 17980
rect 6380 17920 6444 17924
rect 6460 17980 6524 17984
rect 6460 17924 6464 17980
rect 6464 17924 6520 17980
rect 6520 17924 6524 17980
rect 6460 17920 6524 17924
rect 6540 17980 6604 17984
rect 6540 17924 6544 17980
rect 6544 17924 6600 17980
rect 6600 17924 6604 17980
rect 6540 17920 6604 17924
rect 6620 17980 6684 17984
rect 6620 17924 6624 17980
rect 6624 17924 6680 17980
rect 6680 17924 6684 17980
rect 6620 17920 6684 17924
rect 11808 17980 11872 17984
rect 11808 17924 11812 17980
rect 11812 17924 11868 17980
rect 11868 17924 11872 17980
rect 11808 17920 11872 17924
rect 11888 17980 11952 17984
rect 11888 17924 11892 17980
rect 11892 17924 11948 17980
rect 11948 17924 11952 17980
rect 11888 17920 11952 17924
rect 11968 17980 12032 17984
rect 11968 17924 11972 17980
rect 11972 17924 12028 17980
rect 12028 17924 12032 17980
rect 11968 17920 12032 17924
rect 12048 17980 12112 17984
rect 12048 17924 12052 17980
rect 12052 17924 12108 17980
rect 12108 17924 12112 17980
rect 12048 17920 12112 17924
rect 3666 17436 3730 17440
rect 3666 17380 3670 17436
rect 3670 17380 3726 17436
rect 3726 17380 3730 17436
rect 3666 17376 3730 17380
rect 3746 17436 3810 17440
rect 3746 17380 3750 17436
rect 3750 17380 3806 17436
rect 3806 17380 3810 17436
rect 3746 17376 3810 17380
rect 3826 17436 3890 17440
rect 3826 17380 3830 17436
rect 3830 17380 3886 17436
rect 3886 17380 3890 17436
rect 3826 17376 3890 17380
rect 3906 17436 3970 17440
rect 3906 17380 3910 17436
rect 3910 17380 3966 17436
rect 3966 17380 3970 17436
rect 3906 17376 3970 17380
rect 9094 17436 9158 17440
rect 9094 17380 9098 17436
rect 9098 17380 9154 17436
rect 9154 17380 9158 17436
rect 9094 17376 9158 17380
rect 9174 17436 9238 17440
rect 9174 17380 9178 17436
rect 9178 17380 9234 17436
rect 9234 17380 9238 17436
rect 9174 17376 9238 17380
rect 9254 17436 9318 17440
rect 9254 17380 9258 17436
rect 9258 17380 9314 17436
rect 9314 17380 9318 17436
rect 9254 17376 9318 17380
rect 9334 17436 9398 17440
rect 9334 17380 9338 17436
rect 9338 17380 9394 17436
rect 9394 17380 9398 17436
rect 9334 17376 9398 17380
rect 14522 17436 14586 17440
rect 14522 17380 14526 17436
rect 14526 17380 14582 17436
rect 14582 17380 14586 17436
rect 14522 17376 14586 17380
rect 14602 17436 14666 17440
rect 14602 17380 14606 17436
rect 14606 17380 14662 17436
rect 14662 17380 14666 17436
rect 14602 17376 14666 17380
rect 14682 17436 14746 17440
rect 14682 17380 14686 17436
rect 14686 17380 14742 17436
rect 14742 17380 14746 17436
rect 14682 17376 14746 17380
rect 14762 17436 14826 17440
rect 14762 17380 14766 17436
rect 14766 17380 14822 17436
rect 14822 17380 14826 17436
rect 14762 17376 14826 17380
rect 6380 16892 6444 16896
rect 6380 16836 6384 16892
rect 6384 16836 6440 16892
rect 6440 16836 6444 16892
rect 6380 16832 6444 16836
rect 6460 16892 6524 16896
rect 6460 16836 6464 16892
rect 6464 16836 6520 16892
rect 6520 16836 6524 16892
rect 6460 16832 6524 16836
rect 6540 16892 6604 16896
rect 6540 16836 6544 16892
rect 6544 16836 6600 16892
rect 6600 16836 6604 16892
rect 6540 16832 6604 16836
rect 6620 16892 6684 16896
rect 6620 16836 6624 16892
rect 6624 16836 6680 16892
rect 6680 16836 6684 16892
rect 6620 16832 6684 16836
rect 11808 16892 11872 16896
rect 11808 16836 11812 16892
rect 11812 16836 11868 16892
rect 11868 16836 11872 16892
rect 11808 16832 11872 16836
rect 11888 16892 11952 16896
rect 11888 16836 11892 16892
rect 11892 16836 11948 16892
rect 11948 16836 11952 16892
rect 11888 16832 11952 16836
rect 11968 16892 12032 16896
rect 11968 16836 11972 16892
rect 11972 16836 12028 16892
rect 12028 16836 12032 16892
rect 11968 16832 12032 16836
rect 12048 16892 12112 16896
rect 12048 16836 12052 16892
rect 12052 16836 12108 16892
rect 12108 16836 12112 16892
rect 12048 16832 12112 16836
rect 3666 16348 3730 16352
rect 3666 16292 3670 16348
rect 3670 16292 3726 16348
rect 3726 16292 3730 16348
rect 3666 16288 3730 16292
rect 3746 16348 3810 16352
rect 3746 16292 3750 16348
rect 3750 16292 3806 16348
rect 3806 16292 3810 16348
rect 3746 16288 3810 16292
rect 3826 16348 3890 16352
rect 3826 16292 3830 16348
rect 3830 16292 3886 16348
rect 3886 16292 3890 16348
rect 3826 16288 3890 16292
rect 3906 16348 3970 16352
rect 3906 16292 3910 16348
rect 3910 16292 3966 16348
rect 3966 16292 3970 16348
rect 3906 16288 3970 16292
rect 9094 16348 9158 16352
rect 9094 16292 9098 16348
rect 9098 16292 9154 16348
rect 9154 16292 9158 16348
rect 9094 16288 9158 16292
rect 9174 16348 9238 16352
rect 9174 16292 9178 16348
rect 9178 16292 9234 16348
rect 9234 16292 9238 16348
rect 9174 16288 9238 16292
rect 9254 16348 9318 16352
rect 9254 16292 9258 16348
rect 9258 16292 9314 16348
rect 9314 16292 9318 16348
rect 9254 16288 9318 16292
rect 9334 16348 9398 16352
rect 9334 16292 9338 16348
rect 9338 16292 9394 16348
rect 9394 16292 9398 16348
rect 9334 16288 9398 16292
rect 14522 16348 14586 16352
rect 14522 16292 14526 16348
rect 14526 16292 14582 16348
rect 14582 16292 14586 16348
rect 14522 16288 14586 16292
rect 14602 16348 14666 16352
rect 14602 16292 14606 16348
rect 14606 16292 14662 16348
rect 14662 16292 14666 16348
rect 14602 16288 14666 16292
rect 14682 16348 14746 16352
rect 14682 16292 14686 16348
rect 14686 16292 14742 16348
rect 14742 16292 14746 16348
rect 14682 16288 14746 16292
rect 14762 16348 14826 16352
rect 14762 16292 14766 16348
rect 14766 16292 14822 16348
rect 14822 16292 14826 16348
rect 14762 16288 14826 16292
rect 6380 15804 6444 15808
rect 6380 15748 6384 15804
rect 6384 15748 6440 15804
rect 6440 15748 6444 15804
rect 6380 15744 6444 15748
rect 6460 15804 6524 15808
rect 6460 15748 6464 15804
rect 6464 15748 6520 15804
rect 6520 15748 6524 15804
rect 6460 15744 6524 15748
rect 6540 15804 6604 15808
rect 6540 15748 6544 15804
rect 6544 15748 6600 15804
rect 6600 15748 6604 15804
rect 6540 15744 6604 15748
rect 6620 15804 6684 15808
rect 6620 15748 6624 15804
rect 6624 15748 6680 15804
rect 6680 15748 6684 15804
rect 6620 15744 6684 15748
rect 11808 15804 11872 15808
rect 11808 15748 11812 15804
rect 11812 15748 11868 15804
rect 11868 15748 11872 15804
rect 11808 15744 11872 15748
rect 11888 15804 11952 15808
rect 11888 15748 11892 15804
rect 11892 15748 11948 15804
rect 11948 15748 11952 15804
rect 11888 15744 11952 15748
rect 11968 15804 12032 15808
rect 11968 15748 11972 15804
rect 11972 15748 12028 15804
rect 12028 15748 12032 15804
rect 11968 15744 12032 15748
rect 12048 15804 12112 15808
rect 12048 15748 12052 15804
rect 12052 15748 12108 15804
rect 12108 15748 12112 15804
rect 12048 15744 12112 15748
rect 3666 15260 3730 15264
rect 3666 15204 3670 15260
rect 3670 15204 3726 15260
rect 3726 15204 3730 15260
rect 3666 15200 3730 15204
rect 3746 15260 3810 15264
rect 3746 15204 3750 15260
rect 3750 15204 3806 15260
rect 3806 15204 3810 15260
rect 3746 15200 3810 15204
rect 3826 15260 3890 15264
rect 3826 15204 3830 15260
rect 3830 15204 3886 15260
rect 3886 15204 3890 15260
rect 3826 15200 3890 15204
rect 3906 15260 3970 15264
rect 3906 15204 3910 15260
rect 3910 15204 3966 15260
rect 3966 15204 3970 15260
rect 3906 15200 3970 15204
rect 9094 15260 9158 15264
rect 9094 15204 9098 15260
rect 9098 15204 9154 15260
rect 9154 15204 9158 15260
rect 9094 15200 9158 15204
rect 9174 15260 9238 15264
rect 9174 15204 9178 15260
rect 9178 15204 9234 15260
rect 9234 15204 9238 15260
rect 9174 15200 9238 15204
rect 9254 15260 9318 15264
rect 9254 15204 9258 15260
rect 9258 15204 9314 15260
rect 9314 15204 9318 15260
rect 9254 15200 9318 15204
rect 9334 15260 9398 15264
rect 9334 15204 9338 15260
rect 9338 15204 9394 15260
rect 9394 15204 9398 15260
rect 9334 15200 9398 15204
rect 14522 15260 14586 15264
rect 14522 15204 14526 15260
rect 14526 15204 14582 15260
rect 14582 15204 14586 15260
rect 14522 15200 14586 15204
rect 14602 15260 14666 15264
rect 14602 15204 14606 15260
rect 14606 15204 14662 15260
rect 14662 15204 14666 15260
rect 14602 15200 14666 15204
rect 14682 15260 14746 15264
rect 14682 15204 14686 15260
rect 14686 15204 14742 15260
rect 14742 15204 14746 15260
rect 14682 15200 14746 15204
rect 14762 15260 14826 15264
rect 14762 15204 14766 15260
rect 14766 15204 14822 15260
rect 14822 15204 14826 15260
rect 14762 15200 14826 15204
rect 6380 14716 6444 14720
rect 6380 14660 6384 14716
rect 6384 14660 6440 14716
rect 6440 14660 6444 14716
rect 6380 14656 6444 14660
rect 6460 14716 6524 14720
rect 6460 14660 6464 14716
rect 6464 14660 6520 14716
rect 6520 14660 6524 14716
rect 6460 14656 6524 14660
rect 6540 14716 6604 14720
rect 6540 14660 6544 14716
rect 6544 14660 6600 14716
rect 6600 14660 6604 14716
rect 6540 14656 6604 14660
rect 6620 14716 6684 14720
rect 6620 14660 6624 14716
rect 6624 14660 6680 14716
rect 6680 14660 6684 14716
rect 6620 14656 6684 14660
rect 11808 14716 11872 14720
rect 11808 14660 11812 14716
rect 11812 14660 11868 14716
rect 11868 14660 11872 14716
rect 11808 14656 11872 14660
rect 11888 14716 11952 14720
rect 11888 14660 11892 14716
rect 11892 14660 11948 14716
rect 11948 14660 11952 14716
rect 11888 14656 11952 14660
rect 11968 14716 12032 14720
rect 11968 14660 11972 14716
rect 11972 14660 12028 14716
rect 12028 14660 12032 14716
rect 11968 14656 12032 14660
rect 12048 14716 12112 14720
rect 12048 14660 12052 14716
rect 12052 14660 12108 14716
rect 12108 14660 12112 14716
rect 12048 14656 12112 14660
rect 3666 14172 3730 14176
rect 3666 14116 3670 14172
rect 3670 14116 3726 14172
rect 3726 14116 3730 14172
rect 3666 14112 3730 14116
rect 3746 14172 3810 14176
rect 3746 14116 3750 14172
rect 3750 14116 3806 14172
rect 3806 14116 3810 14172
rect 3746 14112 3810 14116
rect 3826 14172 3890 14176
rect 3826 14116 3830 14172
rect 3830 14116 3886 14172
rect 3886 14116 3890 14172
rect 3826 14112 3890 14116
rect 3906 14172 3970 14176
rect 3906 14116 3910 14172
rect 3910 14116 3966 14172
rect 3966 14116 3970 14172
rect 3906 14112 3970 14116
rect 9094 14172 9158 14176
rect 9094 14116 9098 14172
rect 9098 14116 9154 14172
rect 9154 14116 9158 14172
rect 9094 14112 9158 14116
rect 9174 14172 9238 14176
rect 9174 14116 9178 14172
rect 9178 14116 9234 14172
rect 9234 14116 9238 14172
rect 9174 14112 9238 14116
rect 9254 14172 9318 14176
rect 9254 14116 9258 14172
rect 9258 14116 9314 14172
rect 9314 14116 9318 14172
rect 9254 14112 9318 14116
rect 9334 14172 9398 14176
rect 9334 14116 9338 14172
rect 9338 14116 9394 14172
rect 9394 14116 9398 14172
rect 9334 14112 9398 14116
rect 14522 14172 14586 14176
rect 14522 14116 14526 14172
rect 14526 14116 14582 14172
rect 14582 14116 14586 14172
rect 14522 14112 14586 14116
rect 14602 14172 14666 14176
rect 14602 14116 14606 14172
rect 14606 14116 14662 14172
rect 14662 14116 14666 14172
rect 14602 14112 14666 14116
rect 14682 14172 14746 14176
rect 14682 14116 14686 14172
rect 14686 14116 14742 14172
rect 14742 14116 14746 14172
rect 14682 14112 14746 14116
rect 14762 14172 14826 14176
rect 14762 14116 14766 14172
rect 14766 14116 14822 14172
rect 14822 14116 14826 14172
rect 14762 14112 14826 14116
rect 6380 13628 6444 13632
rect 6380 13572 6384 13628
rect 6384 13572 6440 13628
rect 6440 13572 6444 13628
rect 6380 13568 6444 13572
rect 6460 13628 6524 13632
rect 6460 13572 6464 13628
rect 6464 13572 6520 13628
rect 6520 13572 6524 13628
rect 6460 13568 6524 13572
rect 6540 13628 6604 13632
rect 6540 13572 6544 13628
rect 6544 13572 6600 13628
rect 6600 13572 6604 13628
rect 6540 13568 6604 13572
rect 6620 13628 6684 13632
rect 6620 13572 6624 13628
rect 6624 13572 6680 13628
rect 6680 13572 6684 13628
rect 6620 13568 6684 13572
rect 11808 13628 11872 13632
rect 11808 13572 11812 13628
rect 11812 13572 11868 13628
rect 11868 13572 11872 13628
rect 11808 13568 11872 13572
rect 11888 13628 11952 13632
rect 11888 13572 11892 13628
rect 11892 13572 11948 13628
rect 11948 13572 11952 13628
rect 11888 13568 11952 13572
rect 11968 13628 12032 13632
rect 11968 13572 11972 13628
rect 11972 13572 12028 13628
rect 12028 13572 12032 13628
rect 11968 13568 12032 13572
rect 12048 13628 12112 13632
rect 12048 13572 12052 13628
rect 12052 13572 12108 13628
rect 12108 13572 12112 13628
rect 12048 13568 12112 13572
rect 3666 13084 3730 13088
rect 3666 13028 3670 13084
rect 3670 13028 3726 13084
rect 3726 13028 3730 13084
rect 3666 13024 3730 13028
rect 3746 13084 3810 13088
rect 3746 13028 3750 13084
rect 3750 13028 3806 13084
rect 3806 13028 3810 13084
rect 3746 13024 3810 13028
rect 3826 13084 3890 13088
rect 3826 13028 3830 13084
rect 3830 13028 3886 13084
rect 3886 13028 3890 13084
rect 3826 13024 3890 13028
rect 3906 13084 3970 13088
rect 3906 13028 3910 13084
rect 3910 13028 3966 13084
rect 3966 13028 3970 13084
rect 3906 13024 3970 13028
rect 9094 13084 9158 13088
rect 9094 13028 9098 13084
rect 9098 13028 9154 13084
rect 9154 13028 9158 13084
rect 9094 13024 9158 13028
rect 9174 13084 9238 13088
rect 9174 13028 9178 13084
rect 9178 13028 9234 13084
rect 9234 13028 9238 13084
rect 9174 13024 9238 13028
rect 9254 13084 9318 13088
rect 9254 13028 9258 13084
rect 9258 13028 9314 13084
rect 9314 13028 9318 13084
rect 9254 13024 9318 13028
rect 9334 13084 9398 13088
rect 9334 13028 9338 13084
rect 9338 13028 9394 13084
rect 9394 13028 9398 13084
rect 9334 13024 9398 13028
rect 14522 13084 14586 13088
rect 14522 13028 14526 13084
rect 14526 13028 14582 13084
rect 14582 13028 14586 13084
rect 14522 13024 14586 13028
rect 14602 13084 14666 13088
rect 14602 13028 14606 13084
rect 14606 13028 14662 13084
rect 14662 13028 14666 13084
rect 14602 13024 14666 13028
rect 14682 13084 14746 13088
rect 14682 13028 14686 13084
rect 14686 13028 14742 13084
rect 14742 13028 14746 13084
rect 14682 13024 14746 13028
rect 14762 13084 14826 13088
rect 14762 13028 14766 13084
rect 14766 13028 14822 13084
rect 14822 13028 14826 13084
rect 14762 13024 14826 13028
rect 6380 12540 6444 12544
rect 6380 12484 6384 12540
rect 6384 12484 6440 12540
rect 6440 12484 6444 12540
rect 6380 12480 6444 12484
rect 6460 12540 6524 12544
rect 6460 12484 6464 12540
rect 6464 12484 6520 12540
rect 6520 12484 6524 12540
rect 6460 12480 6524 12484
rect 6540 12540 6604 12544
rect 6540 12484 6544 12540
rect 6544 12484 6600 12540
rect 6600 12484 6604 12540
rect 6540 12480 6604 12484
rect 6620 12540 6684 12544
rect 6620 12484 6624 12540
rect 6624 12484 6680 12540
rect 6680 12484 6684 12540
rect 6620 12480 6684 12484
rect 11808 12540 11872 12544
rect 11808 12484 11812 12540
rect 11812 12484 11868 12540
rect 11868 12484 11872 12540
rect 11808 12480 11872 12484
rect 11888 12540 11952 12544
rect 11888 12484 11892 12540
rect 11892 12484 11948 12540
rect 11948 12484 11952 12540
rect 11888 12480 11952 12484
rect 11968 12540 12032 12544
rect 11968 12484 11972 12540
rect 11972 12484 12028 12540
rect 12028 12484 12032 12540
rect 11968 12480 12032 12484
rect 12048 12540 12112 12544
rect 12048 12484 12052 12540
rect 12052 12484 12108 12540
rect 12108 12484 12112 12540
rect 12048 12480 12112 12484
rect 3666 11996 3730 12000
rect 3666 11940 3670 11996
rect 3670 11940 3726 11996
rect 3726 11940 3730 11996
rect 3666 11936 3730 11940
rect 3746 11996 3810 12000
rect 3746 11940 3750 11996
rect 3750 11940 3806 11996
rect 3806 11940 3810 11996
rect 3746 11936 3810 11940
rect 3826 11996 3890 12000
rect 3826 11940 3830 11996
rect 3830 11940 3886 11996
rect 3886 11940 3890 11996
rect 3826 11936 3890 11940
rect 3906 11996 3970 12000
rect 3906 11940 3910 11996
rect 3910 11940 3966 11996
rect 3966 11940 3970 11996
rect 3906 11936 3970 11940
rect 9094 11996 9158 12000
rect 9094 11940 9098 11996
rect 9098 11940 9154 11996
rect 9154 11940 9158 11996
rect 9094 11936 9158 11940
rect 9174 11996 9238 12000
rect 9174 11940 9178 11996
rect 9178 11940 9234 11996
rect 9234 11940 9238 11996
rect 9174 11936 9238 11940
rect 9254 11996 9318 12000
rect 9254 11940 9258 11996
rect 9258 11940 9314 11996
rect 9314 11940 9318 11996
rect 9254 11936 9318 11940
rect 9334 11996 9398 12000
rect 9334 11940 9338 11996
rect 9338 11940 9394 11996
rect 9394 11940 9398 11996
rect 9334 11936 9398 11940
rect 14522 11996 14586 12000
rect 14522 11940 14526 11996
rect 14526 11940 14582 11996
rect 14582 11940 14586 11996
rect 14522 11936 14586 11940
rect 14602 11996 14666 12000
rect 14602 11940 14606 11996
rect 14606 11940 14662 11996
rect 14662 11940 14666 11996
rect 14602 11936 14666 11940
rect 14682 11996 14746 12000
rect 14682 11940 14686 11996
rect 14686 11940 14742 11996
rect 14742 11940 14746 11996
rect 14682 11936 14746 11940
rect 14762 11996 14826 12000
rect 14762 11940 14766 11996
rect 14766 11940 14822 11996
rect 14822 11940 14826 11996
rect 14762 11936 14826 11940
rect 6380 11452 6444 11456
rect 6380 11396 6384 11452
rect 6384 11396 6440 11452
rect 6440 11396 6444 11452
rect 6380 11392 6444 11396
rect 6460 11452 6524 11456
rect 6460 11396 6464 11452
rect 6464 11396 6520 11452
rect 6520 11396 6524 11452
rect 6460 11392 6524 11396
rect 6540 11452 6604 11456
rect 6540 11396 6544 11452
rect 6544 11396 6600 11452
rect 6600 11396 6604 11452
rect 6540 11392 6604 11396
rect 6620 11452 6684 11456
rect 6620 11396 6624 11452
rect 6624 11396 6680 11452
rect 6680 11396 6684 11452
rect 6620 11392 6684 11396
rect 11808 11452 11872 11456
rect 11808 11396 11812 11452
rect 11812 11396 11868 11452
rect 11868 11396 11872 11452
rect 11808 11392 11872 11396
rect 11888 11452 11952 11456
rect 11888 11396 11892 11452
rect 11892 11396 11948 11452
rect 11948 11396 11952 11452
rect 11888 11392 11952 11396
rect 11968 11452 12032 11456
rect 11968 11396 11972 11452
rect 11972 11396 12028 11452
rect 12028 11396 12032 11452
rect 11968 11392 12032 11396
rect 12048 11452 12112 11456
rect 12048 11396 12052 11452
rect 12052 11396 12108 11452
rect 12108 11396 12112 11452
rect 12048 11392 12112 11396
rect 3666 10908 3730 10912
rect 3666 10852 3670 10908
rect 3670 10852 3726 10908
rect 3726 10852 3730 10908
rect 3666 10848 3730 10852
rect 3746 10908 3810 10912
rect 3746 10852 3750 10908
rect 3750 10852 3806 10908
rect 3806 10852 3810 10908
rect 3746 10848 3810 10852
rect 3826 10908 3890 10912
rect 3826 10852 3830 10908
rect 3830 10852 3886 10908
rect 3886 10852 3890 10908
rect 3826 10848 3890 10852
rect 3906 10908 3970 10912
rect 3906 10852 3910 10908
rect 3910 10852 3966 10908
rect 3966 10852 3970 10908
rect 3906 10848 3970 10852
rect 9094 10908 9158 10912
rect 9094 10852 9098 10908
rect 9098 10852 9154 10908
rect 9154 10852 9158 10908
rect 9094 10848 9158 10852
rect 9174 10908 9238 10912
rect 9174 10852 9178 10908
rect 9178 10852 9234 10908
rect 9234 10852 9238 10908
rect 9174 10848 9238 10852
rect 9254 10908 9318 10912
rect 9254 10852 9258 10908
rect 9258 10852 9314 10908
rect 9314 10852 9318 10908
rect 9254 10848 9318 10852
rect 9334 10908 9398 10912
rect 9334 10852 9338 10908
rect 9338 10852 9394 10908
rect 9394 10852 9398 10908
rect 9334 10848 9398 10852
rect 14522 10908 14586 10912
rect 14522 10852 14526 10908
rect 14526 10852 14582 10908
rect 14582 10852 14586 10908
rect 14522 10848 14586 10852
rect 14602 10908 14666 10912
rect 14602 10852 14606 10908
rect 14606 10852 14662 10908
rect 14662 10852 14666 10908
rect 14602 10848 14666 10852
rect 14682 10908 14746 10912
rect 14682 10852 14686 10908
rect 14686 10852 14742 10908
rect 14742 10852 14746 10908
rect 14682 10848 14746 10852
rect 14762 10908 14826 10912
rect 14762 10852 14766 10908
rect 14766 10852 14822 10908
rect 14822 10852 14826 10908
rect 14762 10848 14826 10852
rect 6380 10364 6444 10368
rect 6380 10308 6384 10364
rect 6384 10308 6440 10364
rect 6440 10308 6444 10364
rect 6380 10304 6444 10308
rect 6460 10364 6524 10368
rect 6460 10308 6464 10364
rect 6464 10308 6520 10364
rect 6520 10308 6524 10364
rect 6460 10304 6524 10308
rect 6540 10364 6604 10368
rect 6540 10308 6544 10364
rect 6544 10308 6600 10364
rect 6600 10308 6604 10364
rect 6540 10304 6604 10308
rect 6620 10364 6684 10368
rect 6620 10308 6624 10364
rect 6624 10308 6680 10364
rect 6680 10308 6684 10364
rect 6620 10304 6684 10308
rect 11808 10364 11872 10368
rect 11808 10308 11812 10364
rect 11812 10308 11868 10364
rect 11868 10308 11872 10364
rect 11808 10304 11872 10308
rect 11888 10364 11952 10368
rect 11888 10308 11892 10364
rect 11892 10308 11948 10364
rect 11948 10308 11952 10364
rect 11888 10304 11952 10308
rect 11968 10364 12032 10368
rect 11968 10308 11972 10364
rect 11972 10308 12028 10364
rect 12028 10308 12032 10364
rect 11968 10304 12032 10308
rect 12048 10364 12112 10368
rect 12048 10308 12052 10364
rect 12052 10308 12108 10364
rect 12108 10308 12112 10364
rect 12048 10304 12112 10308
rect 3666 9820 3730 9824
rect 3666 9764 3670 9820
rect 3670 9764 3726 9820
rect 3726 9764 3730 9820
rect 3666 9760 3730 9764
rect 3746 9820 3810 9824
rect 3746 9764 3750 9820
rect 3750 9764 3806 9820
rect 3806 9764 3810 9820
rect 3746 9760 3810 9764
rect 3826 9820 3890 9824
rect 3826 9764 3830 9820
rect 3830 9764 3886 9820
rect 3886 9764 3890 9820
rect 3826 9760 3890 9764
rect 3906 9820 3970 9824
rect 3906 9764 3910 9820
rect 3910 9764 3966 9820
rect 3966 9764 3970 9820
rect 3906 9760 3970 9764
rect 9094 9820 9158 9824
rect 9094 9764 9098 9820
rect 9098 9764 9154 9820
rect 9154 9764 9158 9820
rect 9094 9760 9158 9764
rect 9174 9820 9238 9824
rect 9174 9764 9178 9820
rect 9178 9764 9234 9820
rect 9234 9764 9238 9820
rect 9174 9760 9238 9764
rect 9254 9820 9318 9824
rect 9254 9764 9258 9820
rect 9258 9764 9314 9820
rect 9314 9764 9318 9820
rect 9254 9760 9318 9764
rect 9334 9820 9398 9824
rect 9334 9764 9338 9820
rect 9338 9764 9394 9820
rect 9394 9764 9398 9820
rect 9334 9760 9398 9764
rect 14522 9820 14586 9824
rect 14522 9764 14526 9820
rect 14526 9764 14582 9820
rect 14582 9764 14586 9820
rect 14522 9760 14586 9764
rect 14602 9820 14666 9824
rect 14602 9764 14606 9820
rect 14606 9764 14662 9820
rect 14662 9764 14666 9820
rect 14602 9760 14666 9764
rect 14682 9820 14746 9824
rect 14682 9764 14686 9820
rect 14686 9764 14742 9820
rect 14742 9764 14746 9820
rect 14682 9760 14746 9764
rect 14762 9820 14826 9824
rect 14762 9764 14766 9820
rect 14766 9764 14822 9820
rect 14822 9764 14826 9820
rect 14762 9760 14826 9764
rect 6380 9276 6444 9280
rect 6380 9220 6384 9276
rect 6384 9220 6440 9276
rect 6440 9220 6444 9276
rect 6380 9216 6444 9220
rect 6460 9276 6524 9280
rect 6460 9220 6464 9276
rect 6464 9220 6520 9276
rect 6520 9220 6524 9276
rect 6460 9216 6524 9220
rect 6540 9276 6604 9280
rect 6540 9220 6544 9276
rect 6544 9220 6600 9276
rect 6600 9220 6604 9276
rect 6540 9216 6604 9220
rect 6620 9276 6684 9280
rect 6620 9220 6624 9276
rect 6624 9220 6680 9276
rect 6680 9220 6684 9276
rect 6620 9216 6684 9220
rect 11808 9276 11872 9280
rect 11808 9220 11812 9276
rect 11812 9220 11868 9276
rect 11868 9220 11872 9276
rect 11808 9216 11872 9220
rect 11888 9276 11952 9280
rect 11888 9220 11892 9276
rect 11892 9220 11948 9276
rect 11948 9220 11952 9276
rect 11888 9216 11952 9220
rect 11968 9276 12032 9280
rect 11968 9220 11972 9276
rect 11972 9220 12028 9276
rect 12028 9220 12032 9276
rect 11968 9216 12032 9220
rect 12048 9276 12112 9280
rect 12048 9220 12052 9276
rect 12052 9220 12108 9276
rect 12108 9220 12112 9276
rect 12048 9216 12112 9220
rect 3666 8732 3730 8736
rect 3666 8676 3670 8732
rect 3670 8676 3726 8732
rect 3726 8676 3730 8732
rect 3666 8672 3730 8676
rect 3746 8732 3810 8736
rect 3746 8676 3750 8732
rect 3750 8676 3806 8732
rect 3806 8676 3810 8732
rect 3746 8672 3810 8676
rect 3826 8732 3890 8736
rect 3826 8676 3830 8732
rect 3830 8676 3886 8732
rect 3886 8676 3890 8732
rect 3826 8672 3890 8676
rect 3906 8732 3970 8736
rect 3906 8676 3910 8732
rect 3910 8676 3966 8732
rect 3966 8676 3970 8732
rect 3906 8672 3970 8676
rect 9094 8732 9158 8736
rect 9094 8676 9098 8732
rect 9098 8676 9154 8732
rect 9154 8676 9158 8732
rect 9094 8672 9158 8676
rect 9174 8732 9238 8736
rect 9174 8676 9178 8732
rect 9178 8676 9234 8732
rect 9234 8676 9238 8732
rect 9174 8672 9238 8676
rect 9254 8732 9318 8736
rect 9254 8676 9258 8732
rect 9258 8676 9314 8732
rect 9314 8676 9318 8732
rect 9254 8672 9318 8676
rect 9334 8732 9398 8736
rect 9334 8676 9338 8732
rect 9338 8676 9394 8732
rect 9394 8676 9398 8732
rect 9334 8672 9398 8676
rect 14522 8732 14586 8736
rect 14522 8676 14526 8732
rect 14526 8676 14582 8732
rect 14582 8676 14586 8732
rect 14522 8672 14586 8676
rect 14602 8732 14666 8736
rect 14602 8676 14606 8732
rect 14606 8676 14662 8732
rect 14662 8676 14666 8732
rect 14602 8672 14666 8676
rect 14682 8732 14746 8736
rect 14682 8676 14686 8732
rect 14686 8676 14742 8732
rect 14742 8676 14746 8732
rect 14682 8672 14746 8676
rect 14762 8732 14826 8736
rect 14762 8676 14766 8732
rect 14766 8676 14822 8732
rect 14822 8676 14826 8732
rect 14762 8672 14826 8676
rect 6380 8188 6444 8192
rect 6380 8132 6384 8188
rect 6384 8132 6440 8188
rect 6440 8132 6444 8188
rect 6380 8128 6444 8132
rect 6460 8188 6524 8192
rect 6460 8132 6464 8188
rect 6464 8132 6520 8188
rect 6520 8132 6524 8188
rect 6460 8128 6524 8132
rect 6540 8188 6604 8192
rect 6540 8132 6544 8188
rect 6544 8132 6600 8188
rect 6600 8132 6604 8188
rect 6540 8128 6604 8132
rect 6620 8188 6684 8192
rect 6620 8132 6624 8188
rect 6624 8132 6680 8188
rect 6680 8132 6684 8188
rect 6620 8128 6684 8132
rect 11808 8188 11872 8192
rect 11808 8132 11812 8188
rect 11812 8132 11868 8188
rect 11868 8132 11872 8188
rect 11808 8128 11872 8132
rect 11888 8188 11952 8192
rect 11888 8132 11892 8188
rect 11892 8132 11948 8188
rect 11948 8132 11952 8188
rect 11888 8128 11952 8132
rect 11968 8188 12032 8192
rect 11968 8132 11972 8188
rect 11972 8132 12028 8188
rect 12028 8132 12032 8188
rect 11968 8128 12032 8132
rect 12048 8188 12112 8192
rect 12048 8132 12052 8188
rect 12052 8132 12108 8188
rect 12108 8132 12112 8188
rect 12048 8128 12112 8132
rect 3666 7644 3730 7648
rect 3666 7588 3670 7644
rect 3670 7588 3726 7644
rect 3726 7588 3730 7644
rect 3666 7584 3730 7588
rect 3746 7644 3810 7648
rect 3746 7588 3750 7644
rect 3750 7588 3806 7644
rect 3806 7588 3810 7644
rect 3746 7584 3810 7588
rect 3826 7644 3890 7648
rect 3826 7588 3830 7644
rect 3830 7588 3886 7644
rect 3886 7588 3890 7644
rect 3826 7584 3890 7588
rect 3906 7644 3970 7648
rect 3906 7588 3910 7644
rect 3910 7588 3966 7644
rect 3966 7588 3970 7644
rect 3906 7584 3970 7588
rect 9094 7644 9158 7648
rect 9094 7588 9098 7644
rect 9098 7588 9154 7644
rect 9154 7588 9158 7644
rect 9094 7584 9158 7588
rect 9174 7644 9238 7648
rect 9174 7588 9178 7644
rect 9178 7588 9234 7644
rect 9234 7588 9238 7644
rect 9174 7584 9238 7588
rect 9254 7644 9318 7648
rect 9254 7588 9258 7644
rect 9258 7588 9314 7644
rect 9314 7588 9318 7644
rect 9254 7584 9318 7588
rect 9334 7644 9398 7648
rect 9334 7588 9338 7644
rect 9338 7588 9394 7644
rect 9394 7588 9398 7644
rect 9334 7584 9398 7588
rect 14522 7644 14586 7648
rect 14522 7588 14526 7644
rect 14526 7588 14582 7644
rect 14582 7588 14586 7644
rect 14522 7584 14586 7588
rect 14602 7644 14666 7648
rect 14602 7588 14606 7644
rect 14606 7588 14662 7644
rect 14662 7588 14666 7644
rect 14602 7584 14666 7588
rect 14682 7644 14746 7648
rect 14682 7588 14686 7644
rect 14686 7588 14742 7644
rect 14742 7588 14746 7644
rect 14682 7584 14746 7588
rect 14762 7644 14826 7648
rect 14762 7588 14766 7644
rect 14766 7588 14822 7644
rect 14822 7588 14826 7644
rect 14762 7584 14826 7588
rect 6380 7100 6444 7104
rect 6380 7044 6384 7100
rect 6384 7044 6440 7100
rect 6440 7044 6444 7100
rect 6380 7040 6444 7044
rect 6460 7100 6524 7104
rect 6460 7044 6464 7100
rect 6464 7044 6520 7100
rect 6520 7044 6524 7100
rect 6460 7040 6524 7044
rect 6540 7100 6604 7104
rect 6540 7044 6544 7100
rect 6544 7044 6600 7100
rect 6600 7044 6604 7100
rect 6540 7040 6604 7044
rect 6620 7100 6684 7104
rect 6620 7044 6624 7100
rect 6624 7044 6680 7100
rect 6680 7044 6684 7100
rect 6620 7040 6684 7044
rect 11808 7100 11872 7104
rect 11808 7044 11812 7100
rect 11812 7044 11868 7100
rect 11868 7044 11872 7100
rect 11808 7040 11872 7044
rect 11888 7100 11952 7104
rect 11888 7044 11892 7100
rect 11892 7044 11948 7100
rect 11948 7044 11952 7100
rect 11888 7040 11952 7044
rect 11968 7100 12032 7104
rect 11968 7044 11972 7100
rect 11972 7044 12028 7100
rect 12028 7044 12032 7100
rect 11968 7040 12032 7044
rect 12048 7100 12112 7104
rect 12048 7044 12052 7100
rect 12052 7044 12108 7100
rect 12108 7044 12112 7100
rect 12048 7040 12112 7044
rect 3666 6556 3730 6560
rect 3666 6500 3670 6556
rect 3670 6500 3726 6556
rect 3726 6500 3730 6556
rect 3666 6496 3730 6500
rect 3746 6556 3810 6560
rect 3746 6500 3750 6556
rect 3750 6500 3806 6556
rect 3806 6500 3810 6556
rect 3746 6496 3810 6500
rect 3826 6556 3890 6560
rect 3826 6500 3830 6556
rect 3830 6500 3886 6556
rect 3886 6500 3890 6556
rect 3826 6496 3890 6500
rect 3906 6556 3970 6560
rect 3906 6500 3910 6556
rect 3910 6500 3966 6556
rect 3966 6500 3970 6556
rect 3906 6496 3970 6500
rect 9094 6556 9158 6560
rect 9094 6500 9098 6556
rect 9098 6500 9154 6556
rect 9154 6500 9158 6556
rect 9094 6496 9158 6500
rect 9174 6556 9238 6560
rect 9174 6500 9178 6556
rect 9178 6500 9234 6556
rect 9234 6500 9238 6556
rect 9174 6496 9238 6500
rect 9254 6556 9318 6560
rect 9254 6500 9258 6556
rect 9258 6500 9314 6556
rect 9314 6500 9318 6556
rect 9254 6496 9318 6500
rect 9334 6556 9398 6560
rect 9334 6500 9338 6556
rect 9338 6500 9394 6556
rect 9394 6500 9398 6556
rect 9334 6496 9398 6500
rect 14522 6556 14586 6560
rect 14522 6500 14526 6556
rect 14526 6500 14582 6556
rect 14582 6500 14586 6556
rect 14522 6496 14586 6500
rect 14602 6556 14666 6560
rect 14602 6500 14606 6556
rect 14606 6500 14662 6556
rect 14662 6500 14666 6556
rect 14602 6496 14666 6500
rect 14682 6556 14746 6560
rect 14682 6500 14686 6556
rect 14686 6500 14742 6556
rect 14742 6500 14746 6556
rect 14682 6496 14746 6500
rect 14762 6556 14826 6560
rect 14762 6500 14766 6556
rect 14766 6500 14822 6556
rect 14822 6500 14826 6556
rect 14762 6496 14826 6500
rect 6380 6012 6444 6016
rect 6380 5956 6384 6012
rect 6384 5956 6440 6012
rect 6440 5956 6444 6012
rect 6380 5952 6444 5956
rect 6460 6012 6524 6016
rect 6460 5956 6464 6012
rect 6464 5956 6520 6012
rect 6520 5956 6524 6012
rect 6460 5952 6524 5956
rect 6540 6012 6604 6016
rect 6540 5956 6544 6012
rect 6544 5956 6600 6012
rect 6600 5956 6604 6012
rect 6540 5952 6604 5956
rect 6620 6012 6684 6016
rect 6620 5956 6624 6012
rect 6624 5956 6680 6012
rect 6680 5956 6684 6012
rect 6620 5952 6684 5956
rect 11808 6012 11872 6016
rect 11808 5956 11812 6012
rect 11812 5956 11868 6012
rect 11868 5956 11872 6012
rect 11808 5952 11872 5956
rect 11888 6012 11952 6016
rect 11888 5956 11892 6012
rect 11892 5956 11948 6012
rect 11948 5956 11952 6012
rect 11888 5952 11952 5956
rect 11968 6012 12032 6016
rect 11968 5956 11972 6012
rect 11972 5956 12028 6012
rect 12028 5956 12032 6012
rect 11968 5952 12032 5956
rect 12048 6012 12112 6016
rect 12048 5956 12052 6012
rect 12052 5956 12108 6012
rect 12108 5956 12112 6012
rect 12048 5952 12112 5956
rect 3666 5468 3730 5472
rect 3666 5412 3670 5468
rect 3670 5412 3726 5468
rect 3726 5412 3730 5468
rect 3666 5408 3730 5412
rect 3746 5468 3810 5472
rect 3746 5412 3750 5468
rect 3750 5412 3806 5468
rect 3806 5412 3810 5468
rect 3746 5408 3810 5412
rect 3826 5468 3890 5472
rect 3826 5412 3830 5468
rect 3830 5412 3886 5468
rect 3886 5412 3890 5468
rect 3826 5408 3890 5412
rect 3906 5468 3970 5472
rect 3906 5412 3910 5468
rect 3910 5412 3966 5468
rect 3966 5412 3970 5468
rect 3906 5408 3970 5412
rect 9094 5468 9158 5472
rect 9094 5412 9098 5468
rect 9098 5412 9154 5468
rect 9154 5412 9158 5468
rect 9094 5408 9158 5412
rect 9174 5468 9238 5472
rect 9174 5412 9178 5468
rect 9178 5412 9234 5468
rect 9234 5412 9238 5468
rect 9174 5408 9238 5412
rect 9254 5468 9318 5472
rect 9254 5412 9258 5468
rect 9258 5412 9314 5468
rect 9314 5412 9318 5468
rect 9254 5408 9318 5412
rect 9334 5468 9398 5472
rect 9334 5412 9338 5468
rect 9338 5412 9394 5468
rect 9394 5412 9398 5468
rect 9334 5408 9398 5412
rect 14522 5468 14586 5472
rect 14522 5412 14526 5468
rect 14526 5412 14582 5468
rect 14582 5412 14586 5468
rect 14522 5408 14586 5412
rect 14602 5468 14666 5472
rect 14602 5412 14606 5468
rect 14606 5412 14662 5468
rect 14662 5412 14666 5468
rect 14602 5408 14666 5412
rect 14682 5468 14746 5472
rect 14682 5412 14686 5468
rect 14686 5412 14742 5468
rect 14742 5412 14746 5468
rect 14682 5408 14746 5412
rect 14762 5468 14826 5472
rect 14762 5412 14766 5468
rect 14766 5412 14822 5468
rect 14822 5412 14826 5468
rect 14762 5408 14826 5412
rect 6380 4924 6444 4928
rect 6380 4868 6384 4924
rect 6384 4868 6440 4924
rect 6440 4868 6444 4924
rect 6380 4864 6444 4868
rect 6460 4924 6524 4928
rect 6460 4868 6464 4924
rect 6464 4868 6520 4924
rect 6520 4868 6524 4924
rect 6460 4864 6524 4868
rect 6540 4924 6604 4928
rect 6540 4868 6544 4924
rect 6544 4868 6600 4924
rect 6600 4868 6604 4924
rect 6540 4864 6604 4868
rect 6620 4924 6684 4928
rect 6620 4868 6624 4924
rect 6624 4868 6680 4924
rect 6680 4868 6684 4924
rect 6620 4864 6684 4868
rect 11808 4924 11872 4928
rect 11808 4868 11812 4924
rect 11812 4868 11868 4924
rect 11868 4868 11872 4924
rect 11808 4864 11872 4868
rect 11888 4924 11952 4928
rect 11888 4868 11892 4924
rect 11892 4868 11948 4924
rect 11948 4868 11952 4924
rect 11888 4864 11952 4868
rect 11968 4924 12032 4928
rect 11968 4868 11972 4924
rect 11972 4868 12028 4924
rect 12028 4868 12032 4924
rect 11968 4864 12032 4868
rect 12048 4924 12112 4928
rect 12048 4868 12052 4924
rect 12052 4868 12108 4924
rect 12108 4868 12112 4924
rect 12048 4864 12112 4868
rect 3666 4380 3730 4384
rect 3666 4324 3670 4380
rect 3670 4324 3726 4380
rect 3726 4324 3730 4380
rect 3666 4320 3730 4324
rect 3746 4380 3810 4384
rect 3746 4324 3750 4380
rect 3750 4324 3806 4380
rect 3806 4324 3810 4380
rect 3746 4320 3810 4324
rect 3826 4380 3890 4384
rect 3826 4324 3830 4380
rect 3830 4324 3886 4380
rect 3886 4324 3890 4380
rect 3826 4320 3890 4324
rect 3906 4380 3970 4384
rect 3906 4324 3910 4380
rect 3910 4324 3966 4380
rect 3966 4324 3970 4380
rect 3906 4320 3970 4324
rect 9094 4380 9158 4384
rect 9094 4324 9098 4380
rect 9098 4324 9154 4380
rect 9154 4324 9158 4380
rect 9094 4320 9158 4324
rect 9174 4380 9238 4384
rect 9174 4324 9178 4380
rect 9178 4324 9234 4380
rect 9234 4324 9238 4380
rect 9174 4320 9238 4324
rect 9254 4380 9318 4384
rect 9254 4324 9258 4380
rect 9258 4324 9314 4380
rect 9314 4324 9318 4380
rect 9254 4320 9318 4324
rect 9334 4380 9398 4384
rect 9334 4324 9338 4380
rect 9338 4324 9394 4380
rect 9394 4324 9398 4380
rect 9334 4320 9398 4324
rect 14522 4380 14586 4384
rect 14522 4324 14526 4380
rect 14526 4324 14582 4380
rect 14582 4324 14586 4380
rect 14522 4320 14586 4324
rect 14602 4380 14666 4384
rect 14602 4324 14606 4380
rect 14606 4324 14662 4380
rect 14662 4324 14666 4380
rect 14602 4320 14666 4324
rect 14682 4380 14746 4384
rect 14682 4324 14686 4380
rect 14686 4324 14742 4380
rect 14742 4324 14746 4380
rect 14682 4320 14746 4324
rect 14762 4380 14826 4384
rect 14762 4324 14766 4380
rect 14766 4324 14822 4380
rect 14822 4324 14826 4380
rect 14762 4320 14826 4324
rect 6380 3836 6444 3840
rect 6380 3780 6384 3836
rect 6384 3780 6440 3836
rect 6440 3780 6444 3836
rect 6380 3776 6444 3780
rect 6460 3836 6524 3840
rect 6460 3780 6464 3836
rect 6464 3780 6520 3836
rect 6520 3780 6524 3836
rect 6460 3776 6524 3780
rect 6540 3836 6604 3840
rect 6540 3780 6544 3836
rect 6544 3780 6600 3836
rect 6600 3780 6604 3836
rect 6540 3776 6604 3780
rect 6620 3836 6684 3840
rect 6620 3780 6624 3836
rect 6624 3780 6680 3836
rect 6680 3780 6684 3836
rect 6620 3776 6684 3780
rect 11808 3836 11872 3840
rect 11808 3780 11812 3836
rect 11812 3780 11868 3836
rect 11868 3780 11872 3836
rect 11808 3776 11872 3780
rect 11888 3836 11952 3840
rect 11888 3780 11892 3836
rect 11892 3780 11948 3836
rect 11948 3780 11952 3836
rect 11888 3776 11952 3780
rect 11968 3836 12032 3840
rect 11968 3780 11972 3836
rect 11972 3780 12028 3836
rect 12028 3780 12032 3836
rect 11968 3776 12032 3780
rect 12048 3836 12112 3840
rect 12048 3780 12052 3836
rect 12052 3780 12108 3836
rect 12108 3780 12112 3836
rect 12048 3776 12112 3780
rect 3666 3292 3730 3296
rect 3666 3236 3670 3292
rect 3670 3236 3726 3292
rect 3726 3236 3730 3292
rect 3666 3232 3730 3236
rect 3746 3292 3810 3296
rect 3746 3236 3750 3292
rect 3750 3236 3806 3292
rect 3806 3236 3810 3292
rect 3746 3232 3810 3236
rect 3826 3292 3890 3296
rect 3826 3236 3830 3292
rect 3830 3236 3886 3292
rect 3886 3236 3890 3292
rect 3826 3232 3890 3236
rect 3906 3292 3970 3296
rect 3906 3236 3910 3292
rect 3910 3236 3966 3292
rect 3966 3236 3970 3292
rect 3906 3232 3970 3236
rect 9094 3292 9158 3296
rect 9094 3236 9098 3292
rect 9098 3236 9154 3292
rect 9154 3236 9158 3292
rect 9094 3232 9158 3236
rect 9174 3292 9238 3296
rect 9174 3236 9178 3292
rect 9178 3236 9234 3292
rect 9234 3236 9238 3292
rect 9174 3232 9238 3236
rect 9254 3292 9318 3296
rect 9254 3236 9258 3292
rect 9258 3236 9314 3292
rect 9314 3236 9318 3292
rect 9254 3232 9318 3236
rect 9334 3292 9398 3296
rect 9334 3236 9338 3292
rect 9338 3236 9394 3292
rect 9394 3236 9398 3292
rect 9334 3232 9398 3236
rect 14522 3292 14586 3296
rect 14522 3236 14526 3292
rect 14526 3236 14582 3292
rect 14582 3236 14586 3292
rect 14522 3232 14586 3236
rect 14602 3292 14666 3296
rect 14602 3236 14606 3292
rect 14606 3236 14662 3292
rect 14662 3236 14666 3292
rect 14602 3232 14666 3236
rect 14682 3292 14746 3296
rect 14682 3236 14686 3292
rect 14686 3236 14742 3292
rect 14742 3236 14746 3292
rect 14682 3232 14746 3236
rect 14762 3292 14826 3296
rect 14762 3236 14766 3292
rect 14766 3236 14822 3292
rect 14822 3236 14826 3292
rect 14762 3232 14826 3236
rect 6380 2748 6444 2752
rect 6380 2692 6384 2748
rect 6384 2692 6440 2748
rect 6440 2692 6444 2748
rect 6380 2688 6444 2692
rect 6460 2748 6524 2752
rect 6460 2692 6464 2748
rect 6464 2692 6520 2748
rect 6520 2692 6524 2748
rect 6460 2688 6524 2692
rect 6540 2748 6604 2752
rect 6540 2692 6544 2748
rect 6544 2692 6600 2748
rect 6600 2692 6604 2748
rect 6540 2688 6604 2692
rect 6620 2748 6684 2752
rect 6620 2692 6624 2748
rect 6624 2692 6680 2748
rect 6680 2692 6684 2748
rect 6620 2688 6684 2692
rect 11808 2748 11872 2752
rect 11808 2692 11812 2748
rect 11812 2692 11868 2748
rect 11868 2692 11872 2748
rect 11808 2688 11872 2692
rect 11888 2748 11952 2752
rect 11888 2692 11892 2748
rect 11892 2692 11948 2748
rect 11948 2692 11952 2748
rect 11888 2688 11952 2692
rect 11968 2748 12032 2752
rect 11968 2692 11972 2748
rect 11972 2692 12028 2748
rect 12028 2692 12032 2748
rect 11968 2688 12032 2692
rect 12048 2748 12112 2752
rect 12048 2692 12052 2748
rect 12052 2692 12108 2748
rect 12108 2692 12112 2748
rect 12048 2688 12112 2692
rect 3666 2204 3730 2208
rect 3666 2148 3670 2204
rect 3670 2148 3726 2204
rect 3726 2148 3730 2204
rect 3666 2144 3730 2148
rect 3746 2204 3810 2208
rect 3746 2148 3750 2204
rect 3750 2148 3806 2204
rect 3806 2148 3810 2204
rect 3746 2144 3810 2148
rect 3826 2204 3890 2208
rect 3826 2148 3830 2204
rect 3830 2148 3886 2204
rect 3886 2148 3890 2204
rect 3826 2144 3890 2148
rect 3906 2204 3970 2208
rect 3906 2148 3910 2204
rect 3910 2148 3966 2204
rect 3966 2148 3970 2204
rect 3906 2144 3970 2148
rect 9094 2204 9158 2208
rect 9094 2148 9098 2204
rect 9098 2148 9154 2204
rect 9154 2148 9158 2204
rect 9094 2144 9158 2148
rect 9174 2204 9238 2208
rect 9174 2148 9178 2204
rect 9178 2148 9234 2204
rect 9234 2148 9238 2204
rect 9174 2144 9238 2148
rect 9254 2204 9318 2208
rect 9254 2148 9258 2204
rect 9258 2148 9314 2204
rect 9314 2148 9318 2204
rect 9254 2144 9318 2148
rect 9334 2204 9398 2208
rect 9334 2148 9338 2204
rect 9338 2148 9394 2204
rect 9394 2148 9398 2204
rect 9334 2144 9398 2148
rect 14522 2204 14586 2208
rect 14522 2148 14526 2204
rect 14526 2148 14582 2204
rect 14582 2148 14586 2204
rect 14522 2144 14586 2148
rect 14602 2204 14666 2208
rect 14602 2148 14606 2204
rect 14606 2148 14662 2204
rect 14662 2148 14666 2204
rect 14602 2144 14666 2148
rect 14682 2204 14746 2208
rect 14682 2148 14686 2204
rect 14686 2148 14742 2204
rect 14742 2148 14746 2204
rect 14682 2144 14746 2148
rect 14762 2204 14826 2208
rect 14762 2148 14766 2204
rect 14766 2148 14822 2204
rect 14822 2148 14826 2204
rect 14762 2144 14826 2148
<< metal4 >>
rect 3658 18528 3978 18544
rect 3658 18464 3666 18528
rect 3730 18464 3746 18528
rect 3810 18464 3826 18528
rect 3890 18464 3906 18528
rect 3970 18464 3978 18528
rect 3658 17440 3978 18464
rect 3658 17376 3666 17440
rect 3730 17376 3746 17440
rect 3810 17376 3826 17440
rect 3890 17376 3906 17440
rect 3970 17376 3978 17440
rect 3658 16352 3978 17376
rect 3658 16288 3666 16352
rect 3730 16288 3746 16352
rect 3810 16288 3826 16352
rect 3890 16288 3906 16352
rect 3970 16288 3978 16352
rect 3658 15846 3978 16288
rect 3658 15610 3700 15846
rect 3936 15610 3978 15846
rect 3658 15264 3978 15610
rect 3658 15200 3666 15264
rect 3730 15200 3746 15264
rect 3810 15200 3826 15264
rect 3890 15200 3906 15264
rect 3970 15200 3978 15264
rect 3658 14176 3978 15200
rect 3658 14112 3666 14176
rect 3730 14112 3746 14176
rect 3810 14112 3826 14176
rect 3890 14112 3906 14176
rect 3970 14112 3978 14176
rect 3658 13088 3978 14112
rect 3658 13024 3666 13088
rect 3730 13024 3746 13088
rect 3810 13024 3826 13088
rect 3890 13024 3906 13088
rect 3970 13024 3978 13088
rect 3658 12000 3978 13024
rect 3658 11936 3666 12000
rect 3730 11936 3746 12000
rect 3810 11936 3826 12000
rect 3890 11936 3906 12000
rect 3970 11936 3978 12000
rect 3658 10912 3978 11936
rect 3658 10848 3666 10912
rect 3730 10848 3746 10912
rect 3810 10848 3826 10912
rect 3890 10848 3906 10912
rect 3970 10848 3978 10912
rect 3658 10406 3978 10848
rect 3658 10170 3700 10406
rect 3936 10170 3978 10406
rect 3658 9824 3978 10170
rect 3658 9760 3666 9824
rect 3730 9760 3746 9824
rect 3810 9760 3826 9824
rect 3890 9760 3906 9824
rect 3970 9760 3978 9824
rect 3658 8736 3978 9760
rect 3658 8672 3666 8736
rect 3730 8672 3746 8736
rect 3810 8672 3826 8736
rect 3890 8672 3906 8736
rect 3970 8672 3978 8736
rect 3658 7648 3978 8672
rect 3658 7584 3666 7648
rect 3730 7584 3746 7648
rect 3810 7584 3826 7648
rect 3890 7584 3906 7648
rect 3970 7584 3978 7648
rect 3658 6560 3978 7584
rect 3658 6496 3666 6560
rect 3730 6496 3746 6560
rect 3810 6496 3826 6560
rect 3890 6496 3906 6560
rect 3970 6496 3978 6560
rect 3658 5472 3978 6496
rect 3658 5408 3666 5472
rect 3730 5408 3746 5472
rect 3810 5408 3826 5472
rect 3890 5408 3906 5472
rect 3970 5408 3978 5472
rect 3658 4966 3978 5408
rect 3658 4730 3700 4966
rect 3936 4730 3978 4966
rect 3658 4384 3978 4730
rect 3658 4320 3666 4384
rect 3730 4320 3746 4384
rect 3810 4320 3826 4384
rect 3890 4320 3906 4384
rect 3970 4320 3978 4384
rect 3658 3296 3978 4320
rect 3658 3232 3666 3296
rect 3730 3232 3746 3296
rect 3810 3232 3826 3296
rect 3890 3232 3906 3296
rect 3970 3232 3978 3296
rect 3658 2208 3978 3232
rect 3658 2144 3666 2208
rect 3730 2144 3746 2208
rect 3810 2144 3826 2208
rect 3890 2144 3906 2208
rect 3970 2144 3978 2208
rect 3658 2128 3978 2144
rect 6372 17984 6692 18544
rect 6372 17920 6380 17984
rect 6444 17920 6460 17984
rect 6524 17920 6540 17984
rect 6604 17920 6620 17984
rect 6684 17920 6692 17984
rect 6372 16896 6692 17920
rect 6372 16832 6380 16896
rect 6444 16832 6460 16896
rect 6524 16832 6540 16896
rect 6604 16832 6620 16896
rect 6684 16832 6692 16896
rect 6372 15808 6692 16832
rect 6372 15744 6380 15808
rect 6444 15744 6460 15808
rect 6524 15744 6540 15808
rect 6604 15744 6620 15808
rect 6684 15744 6692 15808
rect 6372 14720 6692 15744
rect 6372 14656 6380 14720
rect 6444 14656 6460 14720
rect 6524 14656 6540 14720
rect 6604 14656 6620 14720
rect 6684 14656 6692 14720
rect 6372 13632 6692 14656
rect 6372 13568 6380 13632
rect 6444 13568 6460 13632
rect 6524 13568 6540 13632
rect 6604 13568 6620 13632
rect 6684 13568 6692 13632
rect 6372 13126 6692 13568
rect 6372 12890 6414 13126
rect 6650 12890 6692 13126
rect 6372 12544 6692 12890
rect 6372 12480 6380 12544
rect 6444 12480 6460 12544
rect 6524 12480 6540 12544
rect 6604 12480 6620 12544
rect 6684 12480 6692 12544
rect 6372 11456 6692 12480
rect 6372 11392 6380 11456
rect 6444 11392 6460 11456
rect 6524 11392 6540 11456
rect 6604 11392 6620 11456
rect 6684 11392 6692 11456
rect 6372 10368 6692 11392
rect 6372 10304 6380 10368
rect 6444 10304 6460 10368
rect 6524 10304 6540 10368
rect 6604 10304 6620 10368
rect 6684 10304 6692 10368
rect 6372 9280 6692 10304
rect 6372 9216 6380 9280
rect 6444 9216 6460 9280
rect 6524 9216 6540 9280
rect 6604 9216 6620 9280
rect 6684 9216 6692 9280
rect 6372 8192 6692 9216
rect 6372 8128 6380 8192
rect 6444 8128 6460 8192
rect 6524 8128 6540 8192
rect 6604 8128 6620 8192
rect 6684 8128 6692 8192
rect 6372 7686 6692 8128
rect 6372 7450 6414 7686
rect 6650 7450 6692 7686
rect 6372 7104 6692 7450
rect 6372 7040 6380 7104
rect 6444 7040 6460 7104
rect 6524 7040 6540 7104
rect 6604 7040 6620 7104
rect 6684 7040 6692 7104
rect 6372 6016 6692 7040
rect 6372 5952 6380 6016
rect 6444 5952 6460 6016
rect 6524 5952 6540 6016
rect 6604 5952 6620 6016
rect 6684 5952 6692 6016
rect 6372 4928 6692 5952
rect 6372 4864 6380 4928
rect 6444 4864 6460 4928
rect 6524 4864 6540 4928
rect 6604 4864 6620 4928
rect 6684 4864 6692 4928
rect 6372 3840 6692 4864
rect 6372 3776 6380 3840
rect 6444 3776 6460 3840
rect 6524 3776 6540 3840
rect 6604 3776 6620 3840
rect 6684 3776 6692 3840
rect 6372 2752 6692 3776
rect 6372 2688 6380 2752
rect 6444 2688 6460 2752
rect 6524 2688 6540 2752
rect 6604 2688 6620 2752
rect 6684 2688 6692 2752
rect 6372 2128 6692 2688
rect 9086 18528 9406 18544
rect 9086 18464 9094 18528
rect 9158 18464 9174 18528
rect 9238 18464 9254 18528
rect 9318 18464 9334 18528
rect 9398 18464 9406 18528
rect 9086 17440 9406 18464
rect 9086 17376 9094 17440
rect 9158 17376 9174 17440
rect 9238 17376 9254 17440
rect 9318 17376 9334 17440
rect 9398 17376 9406 17440
rect 9086 16352 9406 17376
rect 9086 16288 9094 16352
rect 9158 16288 9174 16352
rect 9238 16288 9254 16352
rect 9318 16288 9334 16352
rect 9398 16288 9406 16352
rect 9086 15846 9406 16288
rect 9086 15610 9128 15846
rect 9364 15610 9406 15846
rect 9086 15264 9406 15610
rect 9086 15200 9094 15264
rect 9158 15200 9174 15264
rect 9238 15200 9254 15264
rect 9318 15200 9334 15264
rect 9398 15200 9406 15264
rect 9086 14176 9406 15200
rect 9086 14112 9094 14176
rect 9158 14112 9174 14176
rect 9238 14112 9254 14176
rect 9318 14112 9334 14176
rect 9398 14112 9406 14176
rect 9086 13088 9406 14112
rect 9086 13024 9094 13088
rect 9158 13024 9174 13088
rect 9238 13024 9254 13088
rect 9318 13024 9334 13088
rect 9398 13024 9406 13088
rect 9086 12000 9406 13024
rect 9086 11936 9094 12000
rect 9158 11936 9174 12000
rect 9238 11936 9254 12000
rect 9318 11936 9334 12000
rect 9398 11936 9406 12000
rect 9086 10912 9406 11936
rect 9086 10848 9094 10912
rect 9158 10848 9174 10912
rect 9238 10848 9254 10912
rect 9318 10848 9334 10912
rect 9398 10848 9406 10912
rect 9086 10406 9406 10848
rect 9086 10170 9128 10406
rect 9364 10170 9406 10406
rect 9086 9824 9406 10170
rect 9086 9760 9094 9824
rect 9158 9760 9174 9824
rect 9238 9760 9254 9824
rect 9318 9760 9334 9824
rect 9398 9760 9406 9824
rect 9086 8736 9406 9760
rect 9086 8672 9094 8736
rect 9158 8672 9174 8736
rect 9238 8672 9254 8736
rect 9318 8672 9334 8736
rect 9398 8672 9406 8736
rect 9086 7648 9406 8672
rect 9086 7584 9094 7648
rect 9158 7584 9174 7648
rect 9238 7584 9254 7648
rect 9318 7584 9334 7648
rect 9398 7584 9406 7648
rect 9086 6560 9406 7584
rect 9086 6496 9094 6560
rect 9158 6496 9174 6560
rect 9238 6496 9254 6560
rect 9318 6496 9334 6560
rect 9398 6496 9406 6560
rect 9086 5472 9406 6496
rect 9086 5408 9094 5472
rect 9158 5408 9174 5472
rect 9238 5408 9254 5472
rect 9318 5408 9334 5472
rect 9398 5408 9406 5472
rect 9086 4966 9406 5408
rect 9086 4730 9128 4966
rect 9364 4730 9406 4966
rect 9086 4384 9406 4730
rect 9086 4320 9094 4384
rect 9158 4320 9174 4384
rect 9238 4320 9254 4384
rect 9318 4320 9334 4384
rect 9398 4320 9406 4384
rect 9086 3296 9406 4320
rect 9086 3232 9094 3296
rect 9158 3232 9174 3296
rect 9238 3232 9254 3296
rect 9318 3232 9334 3296
rect 9398 3232 9406 3296
rect 9086 2208 9406 3232
rect 9086 2144 9094 2208
rect 9158 2144 9174 2208
rect 9238 2144 9254 2208
rect 9318 2144 9334 2208
rect 9398 2144 9406 2208
rect 9086 2128 9406 2144
rect 11800 17984 12120 18544
rect 11800 17920 11808 17984
rect 11872 17920 11888 17984
rect 11952 17920 11968 17984
rect 12032 17920 12048 17984
rect 12112 17920 12120 17984
rect 11800 16896 12120 17920
rect 11800 16832 11808 16896
rect 11872 16832 11888 16896
rect 11952 16832 11968 16896
rect 12032 16832 12048 16896
rect 12112 16832 12120 16896
rect 11800 15808 12120 16832
rect 11800 15744 11808 15808
rect 11872 15744 11888 15808
rect 11952 15744 11968 15808
rect 12032 15744 12048 15808
rect 12112 15744 12120 15808
rect 11800 14720 12120 15744
rect 11800 14656 11808 14720
rect 11872 14656 11888 14720
rect 11952 14656 11968 14720
rect 12032 14656 12048 14720
rect 12112 14656 12120 14720
rect 11800 13632 12120 14656
rect 11800 13568 11808 13632
rect 11872 13568 11888 13632
rect 11952 13568 11968 13632
rect 12032 13568 12048 13632
rect 12112 13568 12120 13632
rect 11800 13126 12120 13568
rect 11800 12890 11842 13126
rect 12078 12890 12120 13126
rect 11800 12544 12120 12890
rect 11800 12480 11808 12544
rect 11872 12480 11888 12544
rect 11952 12480 11968 12544
rect 12032 12480 12048 12544
rect 12112 12480 12120 12544
rect 11800 11456 12120 12480
rect 11800 11392 11808 11456
rect 11872 11392 11888 11456
rect 11952 11392 11968 11456
rect 12032 11392 12048 11456
rect 12112 11392 12120 11456
rect 11800 10368 12120 11392
rect 11800 10304 11808 10368
rect 11872 10304 11888 10368
rect 11952 10304 11968 10368
rect 12032 10304 12048 10368
rect 12112 10304 12120 10368
rect 11800 9280 12120 10304
rect 11800 9216 11808 9280
rect 11872 9216 11888 9280
rect 11952 9216 11968 9280
rect 12032 9216 12048 9280
rect 12112 9216 12120 9280
rect 11800 8192 12120 9216
rect 11800 8128 11808 8192
rect 11872 8128 11888 8192
rect 11952 8128 11968 8192
rect 12032 8128 12048 8192
rect 12112 8128 12120 8192
rect 11800 7686 12120 8128
rect 11800 7450 11842 7686
rect 12078 7450 12120 7686
rect 11800 7104 12120 7450
rect 11800 7040 11808 7104
rect 11872 7040 11888 7104
rect 11952 7040 11968 7104
rect 12032 7040 12048 7104
rect 12112 7040 12120 7104
rect 11800 6016 12120 7040
rect 11800 5952 11808 6016
rect 11872 5952 11888 6016
rect 11952 5952 11968 6016
rect 12032 5952 12048 6016
rect 12112 5952 12120 6016
rect 11800 4928 12120 5952
rect 11800 4864 11808 4928
rect 11872 4864 11888 4928
rect 11952 4864 11968 4928
rect 12032 4864 12048 4928
rect 12112 4864 12120 4928
rect 11800 3840 12120 4864
rect 11800 3776 11808 3840
rect 11872 3776 11888 3840
rect 11952 3776 11968 3840
rect 12032 3776 12048 3840
rect 12112 3776 12120 3840
rect 11800 2752 12120 3776
rect 11800 2688 11808 2752
rect 11872 2688 11888 2752
rect 11952 2688 11968 2752
rect 12032 2688 12048 2752
rect 12112 2688 12120 2752
rect 11800 2128 12120 2688
rect 14514 18528 14834 18544
rect 14514 18464 14522 18528
rect 14586 18464 14602 18528
rect 14666 18464 14682 18528
rect 14746 18464 14762 18528
rect 14826 18464 14834 18528
rect 14514 17440 14834 18464
rect 14514 17376 14522 17440
rect 14586 17376 14602 17440
rect 14666 17376 14682 17440
rect 14746 17376 14762 17440
rect 14826 17376 14834 17440
rect 14514 16352 14834 17376
rect 14514 16288 14522 16352
rect 14586 16288 14602 16352
rect 14666 16288 14682 16352
rect 14746 16288 14762 16352
rect 14826 16288 14834 16352
rect 14514 15846 14834 16288
rect 14514 15610 14556 15846
rect 14792 15610 14834 15846
rect 14514 15264 14834 15610
rect 14514 15200 14522 15264
rect 14586 15200 14602 15264
rect 14666 15200 14682 15264
rect 14746 15200 14762 15264
rect 14826 15200 14834 15264
rect 14514 14176 14834 15200
rect 14514 14112 14522 14176
rect 14586 14112 14602 14176
rect 14666 14112 14682 14176
rect 14746 14112 14762 14176
rect 14826 14112 14834 14176
rect 14514 13088 14834 14112
rect 14514 13024 14522 13088
rect 14586 13024 14602 13088
rect 14666 13024 14682 13088
rect 14746 13024 14762 13088
rect 14826 13024 14834 13088
rect 14514 12000 14834 13024
rect 14514 11936 14522 12000
rect 14586 11936 14602 12000
rect 14666 11936 14682 12000
rect 14746 11936 14762 12000
rect 14826 11936 14834 12000
rect 14514 10912 14834 11936
rect 14514 10848 14522 10912
rect 14586 10848 14602 10912
rect 14666 10848 14682 10912
rect 14746 10848 14762 10912
rect 14826 10848 14834 10912
rect 14514 10406 14834 10848
rect 14514 10170 14556 10406
rect 14792 10170 14834 10406
rect 14514 9824 14834 10170
rect 14514 9760 14522 9824
rect 14586 9760 14602 9824
rect 14666 9760 14682 9824
rect 14746 9760 14762 9824
rect 14826 9760 14834 9824
rect 14514 8736 14834 9760
rect 14514 8672 14522 8736
rect 14586 8672 14602 8736
rect 14666 8672 14682 8736
rect 14746 8672 14762 8736
rect 14826 8672 14834 8736
rect 14514 7648 14834 8672
rect 14514 7584 14522 7648
rect 14586 7584 14602 7648
rect 14666 7584 14682 7648
rect 14746 7584 14762 7648
rect 14826 7584 14834 7648
rect 14514 6560 14834 7584
rect 14514 6496 14522 6560
rect 14586 6496 14602 6560
rect 14666 6496 14682 6560
rect 14746 6496 14762 6560
rect 14826 6496 14834 6560
rect 14514 5472 14834 6496
rect 14514 5408 14522 5472
rect 14586 5408 14602 5472
rect 14666 5408 14682 5472
rect 14746 5408 14762 5472
rect 14826 5408 14834 5472
rect 14514 4966 14834 5408
rect 14514 4730 14556 4966
rect 14792 4730 14834 4966
rect 14514 4384 14834 4730
rect 14514 4320 14522 4384
rect 14586 4320 14602 4384
rect 14666 4320 14682 4384
rect 14746 4320 14762 4384
rect 14826 4320 14834 4384
rect 14514 3296 14834 4320
rect 14514 3232 14522 3296
rect 14586 3232 14602 3296
rect 14666 3232 14682 3296
rect 14746 3232 14762 3296
rect 14826 3232 14834 3296
rect 14514 2208 14834 3232
rect 14514 2144 14522 2208
rect 14586 2144 14602 2208
rect 14666 2144 14682 2208
rect 14746 2144 14762 2208
rect 14826 2144 14834 2208
rect 14514 2128 14834 2144
<< via4 >>
rect 3700 15610 3936 15846
rect 3700 10170 3936 10406
rect 3700 4730 3936 4966
rect 6414 12890 6650 13126
rect 6414 7450 6650 7686
rect 9128 15610 9364 15846
rect 9128 10170 9364 10406
rect 9128 4730 9364 4966
rect 11842 12890 12078 13126
rect 11842 7450 12078 7686
rect 14556 15610 14792 15846
rect 14556 10170 14792 10406
rect 14556 4730 14792 4966
<< metal5 >>
rect 1104 15846 17388 15888
rect 1104 15610 3700 15846
rect 3936 15610 9128 15846
rect 9364 15610 14556 15846
rect 14792 15610 17388 15846
rect 1104 15568 17388 15610
rect 1104 13126 17388 13168
rect 1104 12890 6414 13126
rect 6650 12890 11842 13126
rect 12078 12890 17388 13126
rect 1104 12848 17388 12890
rect 1104 10406 17388 10448
rect 1104 10170 3700 10406
rect 3936 10170 9128 10406
rect 9364 10170 14556 10406
rect 14792 10170 17388 10406
rect 1104 10128 17388 10170
rect 1104 7686 17388 7728
rect 1104 7450 6414 7686
rect 6650 7450 11842 7686
rect 12078 7450 17388 7686
rect 1104 7408 17388 7450
rect 1104 4966 17388 5008
rect 1104 4730 3700 4966
rect 3936 4730 9128 4966
rect 9364 4730 14556 4966
rect 14792 4730 17388 4966
rect 1104 4688 17388 4730
use sky130_fd_sc_hd__decap_3  FILLER_1_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 2024 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 1624855595
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 1840 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform -1 0 2024 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1624855595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624855595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 2208 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _405_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform -1 0 3404 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _495_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 2300 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__o2bb2a_1  _406_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 4508 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _407_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 4232 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25
timestamp 1624855595
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1624855595
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1624855595
transform 1 0 4876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_33
timestamp 1624855595
transform 1 0 4140 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1624855595
transform 1 0 5244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45
timestamp 1624855595
transform 1 0 5244 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _431_
timestamp 1624855595
transform 1 0 5336 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _421_
timestamp 1624855595
transform 1 0 5612 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 6440 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_53
timestamp 1624855595
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1624855595
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1624855595
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1624855595
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1624855595
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _265_
timestamp 1624855595
transform -1 0 8740 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _432_
timestamp 1624855595
transform 1 0 6900 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _498_
timestamp 1624855595
transform -1 0 8832 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70
timestamp 1624855595
transform 1 0 7544 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1624855595
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _413_
timestamp 1624855595
transform 1 0 9660 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _416_
timestamp 1624855595
transform 1 0 10488 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 1624855595
transform -1 0 11040 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1624855595
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1624855595
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1624855595
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98
timestamp 1624855595
transform 1 0 10120 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_84
timestamp 1624855595
transform 1 0 8832 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _414_
timestamp 1624855595
transform 1 0 12052 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _499_
timestamp 1624855595
transform -1 0 14076 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1624855595
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1624855595
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110
timestamp 1624855595
transform 1 0 11224 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1624855595
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_108
timestamp 1624855595
transform 1 0 11040 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1624855595
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _266_
timestamp 1624855595
transform 1 0 13156 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _437_
timestamp 1624855595
transform 1 0 14444 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1624855595
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1624855595
transform 1 0 13800 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1624855595
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 1624855595
transform 1 0 12788 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1624855595
transform 1 0 13432 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1624855595
transform 1 0 14076 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _434_
timestamp 1624855595
transform -1 0 15916 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _436_
timestamp 1624855595
transform 1 0 15548 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146
timestamp 1624855595
transform 1 0 14536 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_154
timestamp 1624855595
transform 1 0 15272 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1624855595
transform 1 0 15916 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_153
timestamp 1624855595
transform 1 0 15180 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_164
timestamp 1624855595
transform 1 0 16192 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624855595
transform -1 0 17388 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624855595
transform -1 0 17388 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1624855595
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform -1 0 16744 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1624855595
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_170
timestamp 1624855595
transform 1 0 16744 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_172
timestamp 1624855595
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_1  _408_
timestamp 1624855595
transform 1 0 2668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624855595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1624855595
transform -1 0 2300 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1624855595
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_9
timestamp 1624855595
transform 1 0 1932 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1624855595
transform 1 0 2300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _433_
timestamp 1624855595
transform 1 0 4784 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1624855595
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_25
timestamp 1624855595
transform 1 0 3404 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_30
timestamp 1624855595
transform 1 0 3864 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_38
timestamp 1624855595
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _507_
timestamp 1624855595
transform -1 0 7728 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1624855595
transform 1 0 5520 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _267_
timestamp 1624855595
transform 1 0 8188 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1624855595
transform 1 0 7728 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_76
timestamp 1624855595
transform 1 0 8096 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_80
timestamp 1624855595
transform 1 0 8464 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _412_
timestamp 1624855595
transform 1 0 9476 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624855595
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1624855595
transform -1 0 10856 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1624855595
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1624855595
transform 1 0 10212 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _415_
timestamp 1624855595
transform 1 0 11408 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1624855595
transform 1 0 12420 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_106
timestamp 1624855595
transform 1 0 10856 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 1624855595
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp 1624855595
transform -1 0 13800 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624855595
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_126
timestamp 1624855595
transform 1 0 12696 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_134
timestamp 1624855595
transform 1 0 13432 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_138
timestamp 1624855595
transform 1 0 13800 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_142
timestamp 1624855595
transform 1 0 14168 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_144
timestamp 1624855595
transform 1 0 14352 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _509_
timestamp 1624855595
transform 1 0 14904 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624855595
transform -1 0 17388 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_170
timestamp 1624855595
transform 1 0 16744 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624855595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp 1624855595
transform 1 0 2484 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp 1624855595
transform -1 0 3496 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _430_
timestamp 1624855595
transform -1 0 5244 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1624855595
transform -1 0 4140 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_26
timestamp 1624855595
transform 1 0 3496 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_33
timestamp 1624855595
transform 1 0 4140 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_39
timestamp 1624855595
transform 1 0 4692 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _255_
timestamp 1624855595
transform 1 0 5612 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624855595
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1624855595
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1624855595
transform 1 0 5244 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1624855595
transform 1 0 5888 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_56
timestamp 1624855595
transform 1 0 6256 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_58
timestamp 1624855595
transform 1 0 6440 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _256_
timestamp 1624855595
transform -1 0 8924 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _268_
timestamp 1624855595
transform -1 0 8280 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_65
timestamp 1624855595
transform 1 0 7084 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_73
timestamp 1624855595
transform 1 0 7820 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1624855595
transform 1 0 8280 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _410_
timestamp 1624855595
transform -1 0 10028 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _411_
timestamp 1624855595
transform 1 0 10396 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1624855595
transform 1 0 8924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_97
timestamp 1624855595
transform 1 0 10028 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _263_
timestamp 1624855595
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624855595
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_108
timestamp 1624855595
transform 1 0 11040 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1624855595
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_122
timestamp 1624855595
transform 1 0 12328 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _510_
timestamp 1624855595
transform -1 0 14536 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1624855595
transform 1 0 16192 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _435_
timestamp 1624855595
transform 1 0 15088 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_146
timestamp 1624855595
transform 1 0 14536 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_160
timestamp 1624855595
transform 1 0 15824 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624855595
transform -1 0 17388 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624855595
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_167
timestamp 1624855595
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1624855595
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _270_
timestamp 1624855595
transform -1 0 3036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624855595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1624855595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp 1624855595
transform 1 0 2484 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _508_
timestamp 1624855595
transform 1 0 4232 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624855595
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_21
timestamp 1624855595
transform 1 0 3036 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_30
timestamp 1624855595
transform 1 0 3864 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_54
timestamp 1624855595
transform 1 0 6072 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_62
timestamp 1624855595
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1624855595
transform 1 0 6992 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform -1 0 8648 0 -1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_4_67
timestamp 1624855595
transform 1 0 7268 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_71
timestamp 1624855595
transform 1 0 7636 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_82
timestamp 1624855595
transform 1 0 8648 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _269_
timestamp 1624855595
transform 1 0 9476 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 1624855595
transform 1 0 10212 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624855595
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1624855595
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1624855595
transform 1 0 9752 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_98
timestamp 1624855595
transform 1 0 10120 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _417_
timestamp 1624855595
transform 1 0 12420 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_4_119
timestamp 1624855595
transform 1 0 12052 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1624855595
transform 1 0 13248 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624855595
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1624855595
transform 1 0 12880 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1624855595
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1624855595
transform 1 0 14352 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1624855595
transform -1 0 14996 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1624855595
transform 1 0 16192 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1624855595
transform 1 0 15548 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_151
timestamp 1624855595
transform 1 0 14996 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_160
timestamp 1624855595
transform 1 0 15824 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624855595
transform -1 0 17388 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_167
timestamp 1624855595
transform 1 0 16468 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_173
timestamp 1624855595
transform 1 0 17020 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 1624855595
transform 1 0 1932 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624855595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1624855595
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _400_
timestamp 1624855595
transform 1 0 4140 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_29
timestamp 1624855595
transform 1 0 3772 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_36
timestamp 1624855595
transform 1 0 4416 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _427_
timestamp 1624855595
transform 1 0 5244 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _428_
timestamp 1624855595
transform -1 0 7452 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624855595
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_44
timestamp 1624855595
transform 1 0 5152 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_53
timestamp 1624855595
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_58
timestamp 1624855595
transform 1 0 6440 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _497_
timestamp 1624855595
transform 1 0 7912 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1624855595
transform 1 0 7452 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_73
timestamp 1624855595
transform 1 0 7820 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _420_
timestamp 1624855595
transform 1 0 10488 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_94
timestamp 1624855595
transform 1 0 9752 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 1624855595
transform 1 0 12052 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624855595
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_110
timestamp 1624855595
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_115
timestamp 1624855595
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 1624855595
transform 1 0 14260 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1624855595
transform 1 0 13892 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_163
timestamp 1624855595
transform 1 0 16100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624855595
transform -1 0 17388 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624855595
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_172
timestamp 1624855595
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 1624855595
transform -1 0 2484 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624855595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624855595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1624855595
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_6
timestamp 1624855595
transform 1 0 1656 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_18
timestamp 1624855595
transform 1 0 2760 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1624855595
transform 1 0 1380 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_11
timestamp 1624855595
transform 1 0 2116 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_15
timestamp 1624855595
transform 1 0 2484 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _273_
timestamp 1624855595
transform 1 0 4232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _493_
timestamp 1624855595
transform -1 0 4968 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624855595
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_26
timestamp 1624855595
transform 1 0 3496 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_30
timestamp 1624855595
transform 1 0 3864 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_37
timestamp 1624855595
transform 1 0 4508 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_21
timestamp 1624855595
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _426_
timestamp 1624855595
transform 1 0 5336 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _505_
timestamp 1624855595
transform -1 0 7728 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624855595
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk
timestamp 1624855595
transform 1 0 5612 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_42
timestamp 1624855595
transform 1 0 4968 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1624855595
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_58
timestamp 1624855595
transform 1 0 6440 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1624855595
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _250_
timestamp 1624855595
transform -1 0 8464 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _259_
timestamp 1624855595
transform 1 0 6900 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _424_
timestamp 1624855595
transform -1 0 8556 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 1624855595
transform 1 0 7728 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_80
timestamp 1624855595
transform 1 0 8464 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_66
timestamp 1624855595
transform 1 0 7176 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1624855595
transform 1 0 8556 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _409_
timestamp 1624855595
transform 1 0 9844 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _504_
timestamp 1624855595
transform 1 0 9016 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624855595
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1624855595
transform 1 0 10672 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_87
timestamp 1624855595
transform 1 0 9108 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_100
timestamp 1624855595
transform 1 0 10304 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_85
timestamp 1624855595
transform 1 0 8924 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _418_
timestamp 1624855595
transform 1 0 11316 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _419_
timestamp 1624855595
transform -1 0 13064 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624855595
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk
timestamp 1624855595
transform -1 0 12328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_107
timestamp 1624855595
transform 1 0 10948 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_119
timestamp 1624855595
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_106
timestamp 1624855595
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_115
timestamp 1624855595
transform 1 0 11684 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_122
timestamp 1624855595
transform 1 0 12328 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1624855595
transform -1 0 13432 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _441_
timestamp 1624855595
transform -1 0 14536 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624855595
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1624855595
transform -1 0 13892 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_130
timestamp 1624855595
transform 1 0 13064 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_139
timestamp 1624855595
transform 1 0 13892 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_144
timestamp 1624855595
transform 1 0 14352 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_130
timestamp 1624855595
transform 1 0 13064 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_134
timestamp 1624855595
transform 1 0 13432 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _439_
timestamp 1624855595
transform 1 0 14904 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _511_
timestamp 1624855595
transform 1 0 14904 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1624855595
transform 1 0 16192 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1624855595
transform 1 0 14536 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_158
timestamp 1624855595
transform 1 0 15640 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624855595
transform -1 0 17388 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624855595
transform -1 0 17388 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624855595
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1624855595
transform 1 0 16744 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_167
timestamp 1624855595
transform 1 0 16468 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_172
timestamp 1624855595
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1624855595
transform 1 0 1380 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624855595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 1624855595
transform 1 0 4508 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624855595
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_23
timestamp 1624855595
transform 1 0 3220 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_30
timestamp 1624855595
transform 1 0 3864 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1624855595
transform 1 0 4416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _503_
timestamp 1624855595
transform 1 0 6716 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_8_57
timestamp 1624855595
transform 1 0 6348 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_81
timestamp 1624855595
transform 1 0 8556 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1624855595
transform -1 0 9752 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1624855595
transform 1 0 10120 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624855595
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1624855595
transform 1 0 8924 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1624855595
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_94
timestamp 1624855595
transform 1 0 9752 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_101
timestamp 1624855595
transform 1 0 10396 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _445_
timestamp 1624855595
transform -1 0 12604 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk
timestamp 1624855595
transform -1 0 11040 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_108
timestamp 1624855595
transform 1 0 11040 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_116
timestamp 1624855595
transform 1 0 11776 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_125
timestamp 1624855595
transform 1 0 12604 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _444_
timestamp 1624855595
transform 1 0 12972 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624855595
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_136
timestamp 1624855595
transform 1 0 13616 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_142
timestamp 1624855595
transform 1 0 14168 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_144
timestamp 1624855595
transform 1 0 14352 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _438_
timestamp 1624855595
transform -1 0 16560 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _440_
timestamp 1624855595
transform 1 0 15088 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_8_159
timestamp 1624855595
transform 1 0 15732 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624855595
transform -1 0 17388 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_168
timestamp 1624855595
transform 1 0 16560 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _404_
timestamp 1624855595
transform 1 0 2024 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624855595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1624855595
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1624855595
transform 1 0 1932 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_18
timestamp 1624855595
transform 1 0 2760 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _402_
timestamp 1624855595
transform 1 0 3128 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _403_
timestamp 1624855595
transform -1 0 4876 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1624855595
transform 1 0 3864 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1624855595
transform 1 0 4876 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _258_
timestamp 1624855595
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _429_
timestamp 1624855595
transform 1 0 5244 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624855595
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1624855595
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_58
timestamp 1624855595
transform 1 0 6440 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _423_
timestamp 1624855595
transform -1 0 8464 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk
timestamp 1624855595
transform 1 0 7452 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_65
timestamp 1624855595
transform 1 0 7084 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_80
timestamp 1624855595
transform 1 0 8464 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _425_
timestamp 1624855595
transform -1 0 9568 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _446_
timestamp 1624855595
transform 1 0 10120 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_9_92
timestamp 1624855595
transform 1 0 9568 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_103
timestamp 1624855595
transform 1 0 10580 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _245_
timestamp 1624855595
transform 1 0 10948 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _442_
timestamp 1624855595
transform 1 0 12052 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624855595
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_110
timestamp 1624855595
transform 1 0 11224 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_115
timestamp 1624855595
transform 1 0 11684 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_124
timestamp 1624855595
transform 1 0 12512 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 1624855595
transform 1 0 12972 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_9_128
timestamp 1624855595
transform 1 0 12880 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _422_
timestamp 1624855595
transform -1 0 16100 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_9_149
timestamp 1624855595
transform 1 0 14812 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_157
timestamp 1624855595
transform 1 0 15548 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_163
timestamp 1624855595
transform 1 0 16100 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624855595
transform -1 0 17388 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624855595
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_172
timestamp 1624855595
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _340_
timestamp 1624855595
transform 1 0 2300 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624855595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1624855595
transform 1 0 1748 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1624855595
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_10
timestamp 1624855595
transform 1 0 2024 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1624855595
transform 1 0 2944 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _401_
timestamp 1624855595
transform -1 0 4692 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624855595
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_28
timestamp 1624855595
transform 1 0 3680 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_30
timestamp 1624855595
transform 1 0 3864 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_39
timestamp 1624855595
transform 1 0 4692 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _450_
timestamp 1624855595
transform 1 0 5060 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_10_48
timestamp 1624855595
transform 1 0 5520 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_60
timestamp 1624855595
transform 1 0 6624 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _244_
timestamp 1624855595
transform -1 0 8372 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_72
timestamp 1624855595
transform 1 0 7728 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_79
timestamp 1624855595
transform 1 0 8372 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _516_
timestamp 1624855595
transform 1 0 9752 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624855595
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1624855595
transform -1 0 9752 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1624855595
transform 1 0 8924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1624855595
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _443_
timestamp 1624855595
transform 1 0 11960 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1624855595
transform 1 0 11592 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1624855595
transform -1 0 13892 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624855595
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_126
timestamp 1624855595
transform 1 0 12696 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_134
timestamp 1624855595
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_139
timestamp 1624855595
transform 1 0 13892 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1624855595
transform 1 0 14352 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _363_
timestamp 1624855595
transform -1 0 16008 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk
timestamp 1624855595
transform -1 0 14996 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_151
timestamp 1624855595
transform 1 0 14996 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_162
timestamp 1624855595
transform 1 0 16008 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_166
timestamp 1624855595
transform 1 0 16376 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624855595
transform -1 0 17388 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1624855595
transform 1 0 16468 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1624855595
transform 1 0 16744 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _338_
timestamp 1624855595
transform -1 0 1932 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _463_
timestamp 1624855595
transform -1 0 4416 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624855595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1624855595
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_9
timestamp 1624855595
transform 1 0 1932 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1624855595
transform 1 0 2484 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _336_
timestamp 1624855595
transform 1 0 4784 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_36
timestamp 1624855595
transform 1 0 4416 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _337_
timestamp 1624855595
transform -1 0 5704 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _452_
timestamp 1624855595
transform 1 0 6808 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624855595
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk
timestamp 1624855595
transform -1 0 6348 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_43
timestamp 1624855595
transform 1 0 5060 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_50
timestamp 1624855595
transform 1 0 5704 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_58
timestamp 1624855595
transform 1 0 6440 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _346_
timestamp 1624855595
transform -1 0 8280 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _354_
timestamp 1624855595
transform 1 0 8648 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1624855595
transform 1 0 7452 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_78
timestamp 1624855595
transform 1 0 8280 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _449_
timestamp 1624855595
transform 1 0 9844 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_87
timestamp 1624855595
transform 1 0 9108 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_103
timestamp 1624855595
transform 1 0 10580 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _358_
timestamp 1624855595
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _454_
timestamp 1624855595
transform 1 0 10948 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624855595
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_110
timestamp 1624855595
transform 1 0 11224 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1624855595
transform 1 0 11684 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_122
timestamp 1624855595
transform 1 0 12328 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _513_
timestamp 1624855595
transform -1 0 14628 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_11_126
timestamp 1624855595
transform 1 0 12696 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _366_
timestamp 1624855595
transform 1 0 15088 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1624855595
transform 1 0 16192 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_147
timestamp 1624855595
transform 1 0 14628 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_151
timestamp 1624855595
transform 1 0 14996 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_160
timestamp 1624855595
transform 1 0 15824 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624855595
transform -1 0 17388 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624855595
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_167
timestamp 1624855595
transform 1 0 16468 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1624855595
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_1  _339_
timestamp 1624855595
transform 1 0 2484 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _341_
timestamp 1624855595
transform 1 0 1380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624855595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1624855595
transform 1 0 2116 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _466_
timestamp 1624855595
transform -1 0 6072 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624855595
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_23
timestamp 1624855595
transform 1 0 3220 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_30
timestamp 1624855595
transform 1 0 3864 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _517_
timestamp 1624855595
transform 1 0 6440 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_12_54
timestamp 1624855595
transform 1 0 6072 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_78
timestamp 1624855595
transform 1 0 8280 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _448_
timestamp 1624855595
transform 1 0 9568 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _515_
timestamp 1624855595
transform 1 0 10580 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624855595
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1624855595
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1624855595
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_99
timestamp 1624855595
transform 1 0 10212 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_123
timestamp 1624855595
transform 1 0 12420 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1624855595
transform -1 0 13892 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _367_
timestamp 1624855595
transform 1 0 12788 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624855595
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_132
timestamp 1624855595
transform 1 0 13248 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_139
timestamp 1624855595
transform 1 0 13892 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_144
timestamp 1624855595
transform 1 0 14352 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _475_
timestamp 1624855595
transform 1 0 14904 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624855595
transform -1 0 17388 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1624855595
transform 1 0 16744 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _464_
timestamp 1624855595
transform 1 0 1380 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624855595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624855595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1624855595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1624855595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1624855595
transform -1 0 4876 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1624855595
transform -1 0 3864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624855595
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_30
timestamp 1624855595
transform 1 0 3864 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_41
timestamp 1624855595
transform 1 0 4876 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_23
timestamp 1624855595
transform 1 0 3220 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1624855595
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_47
timestamp 1624855595
transform 1 0 5428 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_42
timestamp 1624855595
transform 1 0 4968 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_1  _453_
timestamp 1624855595
transform -1 0 5980 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1624855595
transform 1 0 5152 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_54
timestamp 1624855595
transform 1 0 6072 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_58
timestamp 1624855595
transform 1 0 6440 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_53
timestamp 1624855595
transform 1 0 5980 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624855595
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1624855595
transform 1 0 5796 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _451_
timestamp 1624855595
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _349_
timestamp 1624855595
transform 1 0 6808 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _348_
timestamp 1624855595
transform 1 0 7912 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _518_
timestamp 1624855595
transform 1 0 8188 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_13_70
timestamp 1624855595
transform 1 0 7544 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_76
timestamp 1624855595
transform 1 0 8096 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_70
timestamp 1624855595
transform 1 0 7544 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_81
timestamp 1624855595
transform 1 0 8556 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _447_
timestamp 1624855595
transform 1 0 10396 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624855595
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform 1 0 9476 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_13_97
timestamp 1624855595
transform 1 0 10028 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1624855595
transform 1 0 8924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1624855595
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1624855595
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _371_
timestamp 1624855595
transform -1 0 12144 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624855595
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_109
timestamp 1624855595
transform 1 0 11132 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1624855595
transform 1 0 11500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1624855595
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_122
timestamp 1624855595
transform 1 0 12328 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_111
timestamp 1624855595
transform 1 0 11316 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_120
timestamp 1624855595
transform 1 0 12144 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _370_
timestamp 1624855595
transform 1 0 12972 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _478_
timestamp 1624855595
transform 1 0 12972 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624855595
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_128
timestamp 1624855595
transform 1 0 12880 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_128
timestamp 1624855595
transform 1 0 12880 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_137
timestamp 1624855595
transform 1 0 13708 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_144
timestamp 1624855595
transform 1 0 14352 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp 1624855595
transform 1 0 16284 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _364_
timestamp 1624855595
transform -1 0 15916 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _365_
timestamp 1624855595
transform -1 0 15916 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_13_149
timestamp 1624855595
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_161
timestamp 1624855595
transform 1 0 15916 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_152
timestamp 1624855595
transform 1 0 15088 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_161
timestamp 1624855595
transform 1 0 15916 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624855595
transform -1 0 17388 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624855595
transform -1 0 17388 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624855595
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1624855595
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_172
timestamp 1624855595
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_168
timestamp 1624855595
transform 1 0 16560 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _398_
timestamp 1624855595
transform 1 0 2024 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624855595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1624855595
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1624855595
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_17
timestamp 1624855595
transform 1 0 2668 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1624855595
transform 1 0 3036 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _472_
timestamp 1624855595
transform 1 0 3680 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1624855595
transform 1 0 3312 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624855595
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1624855595
transform 1 0 5520 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_56
timestamp 1624855595
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_58
timestamp 1624855595
transform 1 0 6440 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _467_
timestamp 1624855595
transform -1 0 9200 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1624855595
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _356_
timestamp 1624855595
transform 1 0 10304 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _357_
timestamp 1624855595
transform 1 0 9568 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1624855595
transform 1 0 9200 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _301_
timestamp 1624855595
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _480_
timestamp 1624855595
transform 1 0 12052 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624855595
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1624855595
transform 1 0 10948 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1624855595
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _368_
timestamp 1624855595
transform -1 0 14996 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_139
timestamp 1624855595
transform 1 0 13892 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _369_
timestamp 1624855595
transform -1 0 16008 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_15_151
timestamp 1624855595
transform 1 0 14996 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_162
timestamp 1624855595
transform 1 0 16008 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624855595
transform -1 0 17388 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624855595
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_170
timestamp 1624855595
transform 1 0 16744 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_172
timestamp 1624855595
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_1  _397_
timestamp 1624855595
transform 1 0 2116 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624855595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1624855595
transform -1 0 2024 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1624855595
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_10
timestamp 1624855595
transform 1 0 2024 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1624855595
transform 1 0 2852 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1624855595
transform 1 0 4508 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624855595
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1624855595
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_30
timestamp 1624855595
transform 1 0 3864 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1624855595
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_57
timestamp 1624855595
transform 1 0 6348 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp 1624855595
transform 1 0 8372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _347_
timestamp 1624855595
transform 1 0 6900 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_71
timestamp 1624855595
transform 1 0 7636 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_82
timestamp 1624855595
transform 1 0 8648 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _471_
timestamp 1624855595
transform -1 0 11408 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624855595
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1624855595
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1624855595
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _374_
timestamp 1624855595
transform -1 0 12512 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_112
timestamp 1624855595
transform 1 0 11408 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_124
timestamp 1624855595
transform 1 0 12512 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1624855595
transform -1 0 13156 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1624855595
transform -1 0 13892 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624855595
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_131
timestamp 1624855595
transform 1 0 13156 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_135
timestamp 1624855595
transform 1 0 13524 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_139
timestamp 1624855595
transform 1 0 13892 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_144
timestamp 1624855595
transform 1 0 14352 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 1624855595
transform 1 0 14904 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624855595
transform -1 0 17388 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1624855595
transform 1 0 16744 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _491_
timestamp 1624855595
transform 1 0 2300 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624855595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1624855595
transform 1 0 1380 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1624855595
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_1  _353_
timestamp 1624855595
transform -1 0 5244 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_33
timestamp 1624855595
transform 1 0 4140 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624855595
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_45
timestamp 1624855595
transform 1 0 5244 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1624855595
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp 1624855595
transform -1 0 7820 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_73
timestamp 1624855595
transform 1 0 7820 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2a_1  _355_
timestamp 1624855595
transform 1 0 10028 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_85
timestamp 1624855595
transform 1 0 8924 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _373_
timestamp 1624855595
transform 1 0 12052 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624855595
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_105
timestamp 1624855595
transform 1 0 10764 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1624855595
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1624855595
transform 1 0 11684 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 1624855595
transform -1 0 15824 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_17_126
timestamp 1624855595
transform 1 0 12696 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_138
timestamp 1624855595
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _295_
timestamp 1624855595
transform 1 0 16192 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_160
timestamp 1624855595
transform 1 0 15824 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624855595
transform -1 0 17388 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624855595
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_167
timestamp 1624855595
transform 1 0 16468 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1624855595
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_1  _399_
timestamp 1624855595
transform 1 0 1380 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624855595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_11
timestamp 1624855595
transform 1 0 2116 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_19
timestamp 1624855595
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _379_
timestamp 1624855595
transform -1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _469_
timestamp 1624855595
transform 1 0 4508 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624855595
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_25
timestamp 1624855595
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_30
timestamp 1624855595
transform 1 0 3864 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1624855595
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _468_
timestamp 1624855595
transform 1 0 6716 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_18_57
timestamp 1624855595
transform 1 0 6348 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_81
timestamp 1624855595
transform 1 0 8556 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _305_
timestamp 1624855595
transform -1 0 10856 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _344_
timestamp 1624855595
transform 1 0 9476 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624855595
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1624855595
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1624855595
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1624855595
transform 1 0 10120 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _291_
timestamp 1624855595
transform -1 0 11776 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _372_
timestamp 1624855595
transform 1 0 12144 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_106
timestamp 1624855595
transform 1 0 10856 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_112
timestamp 1624855595
transform 1 0 11408 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_116
timestamp 1624855595
transform 1 0 11776 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _297_
timestamp 1624855595
transform 1 0 13616 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624855595
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_128
timestamp 1624855595
transform 1 0 12880 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_139
timestamp 1624855595
transform 1 0 13892 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_144
timestamp 1624855595
transform 1 0 14352 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _361_
timestamp 1624855595
transform 1 0 16008 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _362_
timestamp 1624855595
transform 1 0 14904 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_158
timestamp 1624855595
transform 1 0 15640 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624855595
transform -1 0 17388 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_169
timestamp 1624855595
transform 1 0 16652 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_173
timestamp 1624855595
transform 1 0 17020 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _396_
timestamp 1624855595
transform 1 0 1472 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _492_
timestamp 1624855595
transform 1 0 1380 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624855595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624855595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1624855595
transform 1 0 2300 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1624855595
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_9
timestamp 1624855595
transform 1 0 1932 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_16
timestamp 1624855595
transform 1 0 2576 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_23
timestamp 1624855595
transform 1 0 3220 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1624855595
transform 1 0 3680 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_22
timestamp 1624855595
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624855595
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _350_
timestamp 1624855595
transform 1 0 3220 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_20_30
timestamp 1624855595
transform 1 0 3864 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_35
timestamp 1624855595
transform 1 0 4324 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _352_
timestamp 1624855595
transform -1 0 5244 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1624855595
transform 1 0 4048 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _351_
timestamp 1624855595
transform 1 0 4692 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _303_
timestamp 1624855595
transform 1 0 5888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624855595
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk
timestamp 1624855595
transform 1 0 5796 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_47
timestamp 1624855595
transform 1 0 5428 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_54
timestamp 1624855595
transform 1 0 6072 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1624855595
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_45
timestamp 1624855595
transform 1 0 5244 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_51
timestamp 1624855595
transform 1 0 5796 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_55
timestamp 1624855595
transform 1 0 6164 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_67
timestamp 1624855595
transform 1 0 7268 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_63
timestamp 1624855595
transform 1 0 6900 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_70
timestamp 1624855595
transform 1 0 7544 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk
timestamp 1624855595
transform 1 0 7636 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1624855595
transform -1 0 7268 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_74
timestamp 1624855595
transform 1 0 7912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1624855595
transform 1 0 7820 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _345_
timestamp 1624855595
transform 1 0 8096 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _342_
timestamp 1624855595
transform 1 0 8188 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_20_82
timestamp 1624855595
transform 1 0 8648 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _299_
timestamp 1624855595
transform 1 0 10580 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _343_
timestamp 1624855595
transform 1 0 9476 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1624855595
transform 1 0 9384 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624855595
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_84
timestamp 1624855595
transform 1 0 8832 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1624855595
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99
timestamp 1624855595
transform 1 0 10212 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _474_
timestamp 1624855595
transform -1 0 14260 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _479_
timestamp 1624855595
transform -1 0 13064 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624855595
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk
timestamp 1624855595
transform -1 0 12328 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_110
timestamp 1624855595
transform 1 0 11224 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_115
timestamp 1624855595
transform 1 0 11684 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_122
timestamp 1624855595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_106
timestamp 1624855595
transform 1 0 10856 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _287_
timestamp 1624855595
transform 1 0 13524 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624855595
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_143
timestamp 1624855595
transform 1 0 14260 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_130
timestamp 1624855595
transform 1 0 13064 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_134
timestamp 1624855595
transform 1 0 13432 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_139
timestamp 1624855595
transform 1 0 13892 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1624855595
transform 1 0 14352 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _293_
timestamp 1624855595
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _360_
timestamp 1624855595
transform 1 0 15916 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _473_
timestamp 1624855595
transform 1 0 14628 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_20_151
timestamp 1624855595
transform 1 0 14996 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_159
timestamp 1624855595
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624855595
transform -1 0 17388 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624855595
transform -1 0 17388 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624855595
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_167
timestamp 1624855595
transform 1 0 16468 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_172
timestamp 1624855595
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_169
timestamp 1624855595
transform 1 0 16652 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_173
timestamp 1624855595
transform 1 0 17020 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _275_
timestamp 1624855595
transform 1 0 2668 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624855595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1624855595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 1624855595
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_20
timestamp 1624855595
transform 1 0 2944 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _320_
timestamp 1624855595
transform -1 0 3864 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _328_
timestamp 1624855595
transform 1 0 4232 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_21_30
timestamp 1624855595
transform 1 0 3864 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1624855595
transform 1 0 4692 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _331_
timestamp 1624855595
transform -1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _459_
timestamp 1624855595
transform -1 0 8648 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624855595
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1624855595
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_58
timestamp 1624855595
transform 1 0 6440 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1624855595
transform 1 0 8648 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _274_
timestamp 1624855595
transform 1 0 9016 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp 1624855595
transform -1 0 10120 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp 1624855595
transform 1 0 10488 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_90
timestamp 1624855595
transform 1 0 9384 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_94
timestamp 1624855595
transform 1 0 9752 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1624855595
transform 1 0 10120 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1624855595
transform 1 0 12236 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624855595
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk
timestamp 1624855595
transform -1 0 11408 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_105
timestamp 1624855595
transform 1 0 10764 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1624855595
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_115
timestamp 1624855595
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_124
timestamp 1624855595
transform 1 0 12512 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp 1624855595
transform -1 0 14536 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _378_
timestamp 1624855595
transform 1 0 13064 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_138
timestamp 1624855595
transform 1 0 13800 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_142
timestamp 1624855595
transform 1 0 14168 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1624855595
transform 1 0 16100 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1624855595
transform -1 0 15732 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_146
timestamp 1624855595
transform 1 0 14536 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_154
timestamp 1624855595
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1624855595
transform 1 0 15732 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_166
timestamp 1624855595
transform 1 0 16376 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624855595
transform -1 0 17388 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624855595
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_170
timestamp 1624855595
transform 1 0 16744 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1624855595
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _394_
timestamp 1624855595
transform 1 0 2576 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _395_
timestamp 1624855595
transform -1 0 2208 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624855595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1624855595
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_12
timestamp 1624855595
transform 1 0 2208 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _462_
timestamp 1624855595
transform 1 0 4232 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624855595
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_23
timestamp 1624855595
transform 1 0 3220 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_30
timestamp 1624855595
transform 1 0 3864 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _330_
timestamp 1624855595
transform 1 0 6440 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_22_54
timestamp 1624855595
transform 1 0 6072 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _243_
timestamp 1624855595
transform -1 0 8648 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _249_
timestamp 1624855595
transform 1 0 7544 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_65
timestamp 1624855595
transform 1 0 7084 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_69
timestamp 1624855595
transform 1 0 7452 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_74
timestamp 1624855595
transform 1 0 7912 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_82
timestamp 1624855595
transform 1 0 8648 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1624855595
transform -1 0 9752 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _280_
timestamp 1624855595
transform 1 0 10120 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624855595
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1624855595
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_94
timestamp 1624855595
transform 1 0 9752 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_102
timestamp 1624855595
transform 1 0 10488 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _482_
timestamp 1624855595
transform 1 0 11132 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_22_108
timestamp 1624855595
transform 1 0 11040 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624855595
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1624855595
transform 1 0 13616 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_129
timestamp 1624855595
transform 1 0 12972 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_135
timestamp 1624855595
transform 1 0 13524 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_139
timestamp 1624855595
transform 1 0 13892 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1624855595
transform 1 0 14352 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _359_
timestamp 1624855595
transform 1 0 15916 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _376_
timestamp 1624855595
transform 1 0 14720 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_156
timestamp 1624855595
transform 1 0 15456 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_160
timestamp 1624855595
transform 1 0 15824 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_166
timestamp 1624855595
transform 1 0 16376 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624855595
transform -1 0 17388 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1624855595
transform -1 0 4048 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624855595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1624855595
transform 1 0 1748 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1624855595
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_10
timestamp 1624855595
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _278_
timestamp 1624855595
transform 1 0 4416 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_32
timestamp 1624855595
transform 1 0 4048 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_39
timestamp 1624855595
transform 1 0 4692 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _329_
timestamp 1624855595
transform 1 0 5244 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _460_
timestamp 1624855595
transform 1 0 6808 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624855595
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_53
timestamp 1624855595
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_58
timestamp 1624855595
transform 1 0 6440 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_82
timestamp 1624855595
transform 1 0 8648 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1624855595
transform 1 0 9016 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624855595
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1624855595
transform -1 0 12512 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk
timestamp 1624855595
transform -1 0 11592 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_106
timestamp 1624855595
transform 1 0 10856 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_110
timestamp 1624855595
transform 1 0 11224 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_115
timestamp 1624855595
transform 1 0 11684 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_124
timestamp 1624855595
transform 1 0 12512 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _375_
timestamp 1624855595
transform 1 0 12880 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _481_
timestamp 1624855595
transform 1 0 13800 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_23_133
timestamp 1624855595
transform 1 0 13340 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_137
timestamp 1624855595
transform 1 0 13708 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1624855595
transform 1 0 16192 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_158
timestamp 1624855595
transform 1 0 15640 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624855595
transform -1 0 17388 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624855595
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_167
timestamp 1624855595
transform 1 0 16468 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_172
timestamp 1624855595
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_1  _393_
timestamp 1624855595
transform 1 0 1840 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624855595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1624855595
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1624855595
transform 1 0 1748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_16
timestamp 1624855595
transform 1 0 2576 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1624855595
transform -1 0 4692 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624855595
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1624855595
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_30
timestamp 1624855595
transform 1 0 3864 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_39
timestamp 1624855595
transform 1 0 4692 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1624855595
transform -1 0 6256 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk
timestamp 1624855595
transform -1 0 6900 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_51
timestamp 1624855595
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_56
timestamp 1624855595
transform 1 0 6256 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _311_
timestamp 1624855595
transform -1 0 8188 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 1624855595
transform -1 0 7544 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_63
timestamp 1624855595
transform 1 0 6900 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_70
timestamp 1624855595
transform 1 0 7544 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_77
timestamp 1624855595
transform 1 0 8188 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _390_
timestamp 1624855595
transform 1 0 9844 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624855595
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1624855595
transform 1 0 8924 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_87
timestamp 1624855595
transform 1 0 9108 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1624855595
transform 1 0 10488 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _487_
timestamp 1624855595
transform 1 0 10856 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _281_
timestamp 1624855595
transform 1 0 13064 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624855595
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_126
timestamp 1624855595
transform 1 0 12696 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_133
timestamp 1624855595
transform 1 0 13340 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1624855595
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_144
timestamp 1624855595
transform 1 0 14352 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 1624855595
transform 1 0 14904 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624855595
transform -1 0 17388 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_170
timestamp 1624855595
transform 1 0 16744 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _335_
timestamp 1624855595
transform -1 0 3036 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _392_
timestamp 1624855595
transform 1 0 1472 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624855595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1624855595
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_9
timestamp 1624855595
transform 1 0 1932 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp 1624855595
transform 1 0 4416 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _334_
timestamp 1624855595
transform -1 0 4048 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1624855595
transform 1 0 3036 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1624855595
transform 1 0 4048 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_39
timestamp 1624855595
transform 1 0 4692 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1624855595
transform -1 0 5980 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624855595
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_47
timestamp 1624855595
transform 1 0 5428 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_53
timestamp 1624855595
transform 1 0 5980 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_58
timestamp 1624855595
transform 1 0 6440 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1624855595
transform 1 0 8740 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _322_
timestamp 1624855595
transform 1 0 7636 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1624855595
transform -1 0 7268 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_67
timestamp 1624855595
transform 1 0 7268 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_79
timestamp 1624855595
transform 1 0 8372 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp 1624855595
transform 1 0 9384 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _389_
timestamp 1624855595
transform 1 0 10396 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_86
timestamp 1624855595
transform 1 0 9016 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_93
timestamp 1624855595
transform 1 0 9660 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _386_
timestamp 1624855595
transform 1 0 12052 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624855595
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_109
timestamp 1624855595
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1624855595
transform 1 0 11500 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_115
timestamp 1624855595
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1624855595
transform 1 0 13064 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _377_
timestamp 1624855595
transform 1 0 13892 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_126
timestamp 1624855595
transform 1 0 12696 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_133
timestamp 1624855595
transform 1 0 13340 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp 1624855595
transform -1 0 16192 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1624855595
transform 1 0 15272 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_146
timestamp 1624855595
transform 1 0 14536 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_157
timestamp 1624855595
transform 1 0 15548 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_164
timestamp 1624855595
transform 1 0 16192 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624855595
transform -1 0 17388 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624855595
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_170
timestamp 1624855595
transform 1 0 16744 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1624855595
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1624855595
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624855595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624855595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_20
timestamp 1624855595
transform 1 0 2944 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_16
timestamp 1624855595
transform 1 0 2576 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1624855595
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_15
timestamp 1624855595
transform 1 0 2484 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1624855595
transform -1 0 2576 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _333_
timestamp 1624855595
transform 1 0 2576 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1624855595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _458_
timestamp 1624855595
transform 1 0 4876 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _461_
timestamp 1624855595
transform -1 0 4876 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624855595
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1624855595
transform 1 0 3312 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_28
timestamp 1624855595
transform 1 0 3680 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_30
timestamp 1624855595
transform 1 0 3864 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_38
timestamp 1624855595
transform 1 0 4600 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1624855595
transform 1 0 4876 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _324_
timestamp 1624855595
transform 1 0 6808 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _326_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform -1 0 5704 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624855595
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_61
timestamp 1624855595
transform 1 0 6716 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1624855595
transform 1 0 5704 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_56
timestamp 1624855595
transform 1 0 6256 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1624855595
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _323_
timestamp 1624855595
transform 1 0 7636 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _455_
timestamp 1624855595
transform 1 0 7912 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_26_69
timestamp 1624855595
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1624855595
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_70
timestamp 1624855595
transform 1 0 7544 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _388_
timestamp 1624855595
transform -1 0 10948 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _391_
timestamp 1624855595
transform 1 0 9936 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624855595
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_87
timestamp 1624855595
transform 1 0 9108 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_95
timestamp 1624855595
transform 1 0 9844 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_104
timestamp 1624855595
transform 1 0 10672 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_94
timestamp 1624855595
transform 1 0 9752 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform -1 0 11316 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _385_
timestamp 1624855595
transform 1 0 11868 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _485_
timestamp 1624855595
transform -1 0 14076 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624855595
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_111
timestamp 1624855595
transform 1 0 11316 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1624855595
transform 1 0 12604 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_107
timestamp 1624855595
transform 1 0 10948 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1624855595
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_115
timestamp 1624855595
transform 1 0 11684 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _283_
timestamp 1624855595
transform 1 0 13616 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 1624855595
transform -1 0 13248 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624855595
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_132
timestamp 1624855595
transform 1 0 13248 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_139
timestamp 1624855595
transform 1 0 13892 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_144
timestamp 1624855595
transform 1 0 14352 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_141
timestamp 1624855595
transform 1 0 14076 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1624855595
transform 1 0 15916 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _383_
timestamp 1624855595
transform -1 0 15456 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _483_
timestamp 1624855595
transform 1 0 14628 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_26_156
timestamp 1624855595
transform 1 0 15456 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_160
timestamp 1624855595
transform 1 0 15824 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_164
timestamp 1624855595
transform 1 0 16192 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624855595
transform -1 0 17388 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624855595
transform -1 0 17388 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624855595
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_172
timestamp 1624855595
transform 1 0 16928 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_167
timestamp 1624855595
transform 1 0 16468 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_172
timestamp 1624855595
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__and2_1  _321_
timestamp 1624855595
transform 1 0 2944 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _332_
timestamp 1624855595
transform 1 0 2116 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624855595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1624855595
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_16
timestamp 1624855595
transform 1 0 2576 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _457_
timestamp 1624855595
transform -1 0 6440 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624855595
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_25
timestamp 1624855595
transform 1 0 3404 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_30
timestamp 1624855595
transform 1 0 3864 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _456_
timestamp 1624855595
transform 1 0 6808 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1624855595
transform 1 0 6440 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_82
timestamp 1624855595
transform 1 0 8648 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 1624855595
transform 1 0 9476 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624855595
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_87
timestamp 1624855595
transform 1 0 9108 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _486_
timestamp 1624855595
transform 1 0 12052 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_28_111
timestamp 1624855595
transform 1 0 11316 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624855595
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_139
timestamp 1624855595
transform 1 0 13892 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_144
timestamp 1624855595
transform 1 0 14352 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _381_
timestamp 1624855595
transform 1 0 14904 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_158
timestamp 1624855595
transform 1 0 15640 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_166
timestamp 1624855595
transform 1 0 16376 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624855595
transform -1 0 17388 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1624855595
transform 1 0 16468 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1624855595
transform 1 0 16744 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624855595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1624855595
transform -1 0 2024 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1624855595
transform 1 0 2392 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1624855595
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_10
timestamp 1624855595
transform 1 0 2024 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_17
timestamp 1624855595
transform 1 0 2668 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624855595
transform -1 0 5428 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624855595
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1624855595
transform -1 0 3404 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_21
timestamp 1624855595
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_25
timestamp 1624855595
transform 1 0 3404 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_30
timestamp 1624855595
transform 1 0 3864 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_38
timestamp 1624855595
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1624855595
transform 1 0 5796 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624855595
transform 1 0 6440 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_47
timestamp 1624855595
transform 1 0 5428 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_54
timestamp 1624855595
transform 1 0 6072 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_59
timestamp 1624855595
transform 1 0 6532 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp 1624855595
transform 1 0 7176 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output35
timestamp 1624855595
transform -1 0 8188 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_65
timestamp 1624855595
transform 1 0 7084 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1624855595
transform 1 0 7452 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_77
timestamp 1624855595
transform 1 0 8188 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _380_
timestamp 1624855595
transform 1 0 9660 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624855595
transform 1 0 9108 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_85
timestamp 1624855595
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_88
timestamp 1624855595
transform 1 0 9200 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_92
timestamp 1624855595
transform 1 0 9568 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_98
timestamp 1624855595
transform 1 0 10120 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _384_
timestamp 1624855595
transform 1 0 10948 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _387_
timestamp 1624855595
transform -1 0 12972 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624855595
transform 1 0 11776 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_106
timestamp 1624855595
transform 1 0 10856 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_112
timestamp 1624855595
transform 1 0 11408 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_117
timestamp 1624855595
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624855595
transform 1 0 14444 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1624855595
transform 1 0 13340 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_129
timestamp 1624855595
transform 1 0 12972 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_136
timestamp 1624855595
transform 1 0 13616 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_144
timestamp 1624855595
transform 1 0 14352 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _382_
timestamp 1624855595
transform -1 0 15548 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1624855595
transform 1 0 15916 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_146
timestamp 1624855595
transform 1 0 14536 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_157
timestamp 1624855595
transform 1 0 15548 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_164
timestamp 1624855595
transform 1 0 16192 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624855595
transform -1 0 17388 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_172
timestamp 1624855595
transform 1 0 16928 0 1 17952
box -38 -48 222 592
<< labels >>
rlabel metal3 s 0 2728 800 2848 6 clk
port 0 nsew signal input
rlabel metal2 s 7838 19892 7894 20692 6 p
port 1 nsew signal tristate
rlabel metal2 s 11058 19892 11114 20692 6 rst
port 2 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 x[0]
port 3 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 x[10]
port 4 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 x[11]
port 5 nsew signal input
rlabel metal2 s 12898 19892 12954 20692 6 x[12]
port 6 nsew signal input
rlabel metal2 s 9678 19892 9734 20692 6 x[13]
port 7 nsew signal input
rlabel metal2 s 17958 19892 18014 20692 6 x[14]
port 8 nsew signal input
rlabel metal2 s 16578 19892 16634 20692 6 x[15]
port 9 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 x[16]
port 10 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 x[17]
port 11 nsew signal input
rlabel metal2 s 4158 19892 4214 20692 6 x[18]
port 12 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 x[19]
port 13 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 x[1]
port 14 nsew signal input
rlabel metal3 s 17748 12248 18548 12368 6 x[20]
port 15 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 x[21]
port 16 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 x[22]
port 17 nsew signal input
rlabel metal3 s 17748 9528 18548 9648 6 x[23]
port 18 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 x[24]
port 19 nsew signal input
rlabel metal2 s 478 0 534 800 6 x[25]
port 20 nsew signal input
rlabel metal3 s 17748 2048 18548 2168 6 x[26]
port 21 nsew signal input
rlabel metal3 s 17748 14968 18548 15088 6 x[27]
port 22 nsew signal input
rlabel metal3 s 17748 4768 18548 4888 6 x[28]
port 23 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 x[29]
port 24 nsew signal input
rlabel metal2 s 938 19892 994 20692 6 x[2]
port 25 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 x[30]
port 26 nsew signal input
rlabel metal2 s 5998 19892 6054 20692 6 x[31]
port 27 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 x[3]
port 28 nsew signal input
rlabel metal2 s 14738 19892 14794 20692 6 x[4]
port 29 nsew signal input
rlabel metal3 s 17748 7488 18548 7608 6 x[5]
port 30 nsew signal input
rlabel metal2 s 2318 19892 2374 20692 6 x[6]
port 31 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 x[7]
port 32 nsew signal input
rlabel metal3 s 17748 17688 18548 17808 6 x[8]
port 33 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 x[9]
port 34 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 y
port 35 nsew signal input
rlabel metal4 s 14514 2128 14834 18544 6 VPWR
port 36 nsew power bidirectional
rlabel metal4 s 9086 2128 9406 18544 6 VPWR
port 37 nsew power bidirectional
rlabel metal4 s 3658 2128 3978 18544 6 VPWR
port 38 nsew power bidirectional
rlabel metal5 s 1104 15568 17388 15888 6 VPWR
port 39 nsew power bidirectional
rlabel metal5 s 1104 10128 17388 10448 6 VPWR
port 40 nsew power bidirectional
rlabel metal5 s 1104 4688 17388 5008 6 VPWR
port 41 nsew power bidirectional
rlabel metal4 s 11800 2128 12120 18544 6 VGND
port 42 nsew ground bidirectional
rlabel metal4 s 6372 2128 6692 18544 6 VGND
port 43 nsew ground bidirectional
rlabel metal5 s 1104 12848 17388 13168 6 VGND
port 44 nsew ground bidirectional
rlabel metal5 s 1104 7408 17388 7728 6 VGND
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 18548 20692
<< end >>
