magic
tech sky130A
magscale 1 2
timestamp 1738988170
<< obsli1 >>
rect 1104 2159 17388 18513
<< obsm1 >>
rect 474 2048 18018 18544
<< metal2 >>
rect 938 19892 994 20692
rect 2318 19892 2374 20692
rect 4158 19892 4214 20692
rect 5998 19892 6054 20692
rect 7838 19892 7894 20692
rect 9678 19892 9734 20692
rect 11058 19892 11114 20692
rect 12898 19892 12954 20692
rect 14738 19892 14794 20692
rect 16578 19892 16634 20692
rect 17958 19892 18014 20692
rect 478 0 534 800
rect 1858 0 1914 800
rect 3698 0 3754 800
rect 5538 0 5594 800
rect 7378 0 7434 800
rect 8758 0 8814 800
rect 10598 0 10654 800
rect 12438 0 12494 800
rect 14278 0 14334 800
rect 16118 0 16174 800
rect 17498 0 17554 800
<< obsm2 >>
rect 480 19836 882 19892
rect 1050 19836 2262 19892
rect 2430 19836 4102 19892
rect 4270 19836 5942 19892
rect 6110 19836 7782 19892
rect 7950 19836 9622 19892
rect 9790 19836 11002 19892
rect 11170 19836 12842 19892
rect 13010 19836 14682 19892
rect 14850 19836 16522 19892
rect 16690 19836 17902 19892
rect 480 856 18012 19836
rect 590 800 1802 856
rect 1970 800 3642 856
rect 3810 800 5482 856
rect 5650 800 7322 856
rect 7490 800 8702 856
rect 8870 800 10542 856
rect 10710 800 12382 856
rect 12550 800 14222 856
rect 14390 800 16062 856
rect 16230 800 17442 856
rect 17610 800 18012 856
<< metal3 >>
rect 0 18368 800 18488
rect 17748 17688 18548 17808
rect 0 15648 800 15768
rect 17748 14968 18548 15088
rect 0 12928 800 13048
rect 17748 12248 18548 12368
rect 0 10888 800 11008
rect 17748 9528 18548 9648
rect 0 8168 800 8288
rect 17748 7488 18548 7608
rect 0 5448 800 5568
rect 17748 4768 18548 4888
rect 0 2728 800 2848
rect 17748 2048 18548 2168
<< obsm3 >>
rect 880 18288 17748 18529
rect 800 17888 17748 18288
rect 800 17608 17668 17888
rect 800 15848 17748 17608
rect 880 15568 17748 15848
rect 800 15168 17748 15568
rect 800 14888 17668 15168
rect 800 13128 17748 14888
rect 880 12848 17748 13128
rect 800 12448 17748 12848
rect 800 12168 17668 12448
rect 800 11088 17748 12168
rect 880 10808 17748 11088
rect 800 9728 17748 10808
rect 800 9448 17668 9728
rect 800 8368 17748 9448
rect 880 8088 17748 8368
rect 800 7688 17748 8088
rect 800 7408 17668 7688
rect 800 5648 17748 7408
rect 880 5368 17748 5648
rect 800 4968 17748 5368
rect 800 4688 17668 4968
rect 800 2928 17748 4688
rect 880 2648 17748 2928
rect 800 2248 17748 2648
rect 800 2075 17668 2248
<< metal4 >>
rect 3658 2128 3978 18544
rect 6372 2128 6692 18544
rect 9086 2128 9406 18544
rect 11800 2128 12120 18544
rect 14514 2128 14834 18544
<< metal5 >>
rect 1104 15568 17388 15888
rect 1104 12848 17388 13168
rect 1104 10128 17388 10448
rect 1104 7408 17388 7728
rect 1104 4688 17388 5008
<< labels >>
rlabel metal3 s 0 2728 800 2848 6 clk
port 1 nsew signal input
rlabel metal2 s 7838 19892 7894 20692 6 p
port 2 nsew signal output
rlabel metal2 s 11058 19892 11114 20692 6 rst
port 3 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 x[0]
port 4 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 x[10]
port 5 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 x[11]
port 6 nsew signal input
rlabel metal2 s 12898 19892 12954 20692 6 x[12]
port 7 nsew signal input
rlabel metal2 s 9678 19892 9734 20692 6 x[13]
port 8 nsew signal input
rlabel metal2 s 17958 19892 18014 20692 6 x[14]
port 9 nsew signal input
rlabel metal2 s 16578 19892 16634 20692 6 x[15]
port 10 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 x[16]
port 11 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 x[17]
port 12 nsew signal input
rlabel metal2 s 4158 19892 4214 20692 6 x[18]
port 13 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 x[19]
port 14 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 x[1]
port 15 nsew signal input
rlabel metal3 s 17748 12248 18548 12368 6 x[20]
port 16 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 x[21]
port 17 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 x[22]
port 18 nsew signal input
rlabel metal3 s 17748 9528 18548 9648 6 x[23]
port 19 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 x[24]
port 20 nsew signal input
rlabel metal2 s 478 0 534 800 6 x[25]
port 21 nsew signal input
rlabel metal3 s 17748 2048 18548 2168 6 x[26]
port 22 nsew signal input
rlabel metal3 s 17748 14968 18548 15088 6 x[27]
port 23 nsew signal input
rlabel metal3 s 17748 4768 18548 4888 6 x[28]
port 24 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 x[29]
port 25 nsew signal input
rlabel metal2 s 938 19892 994 20692 6 x[2]
port 26 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 x[30]
port 27 nsew signal input
rlabel metal2 s 5998 19892 6054 20692 6 x[31]
port 28 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 x[3]
port 29 nsew signal input
rlabel metal2 s 14738 19892 14794 20692 6 x[4]
port 30 nsew signal input
rlabel metal3 s 17748 7488 18548 7608 6 x[5]
port 31 nsew signal input
rlabel metal2 s 2318 19892 2374 20692 6 x[6]
port 32 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 x[7]
port 33 nsew signal input
rlabel metal3 s 17748 17688 18548 17808 6 x[8]
port 34 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 x[9]
port 35 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 y
port 36 nsew signal input
rlabel metal4 s 14514 2128 14834 18544 6 VPWR
port 37 nsew power bidirectional
rlabel metal4 s 9086 2128 9406 18544 6 VPWR
port 38 nsew power bidirectional
rlabel metal4 s 3658 2128 3978 18544 6 VPWR
port 39 nsew power bidirectional
rlabel metal5 s 1104 15568 17388 15888 6 VPWR
port 40 nsew power bidirectional
rlabel metal5 s 1104 10128 17388 10448 6 VPWR
port 41 nsew power bidirectional
rlabel metal5 s 1104 4688 17388 5008 6 VPWR
port 42 nsew power bidirectional
rlabel metal4 s 11800 2128 12120 18544 6 VGND
port 43 nsew ground bidirectional
rlabel metal4 s 6372 2128 6692 18544 6 VGND
port 44 nsew ground bidirectional
rlabel metal5 s 1104 12848 17388 13168 6 VGND
port 45 nsew ground bidirectional
rlabel metal5 s 1104 7408 17388 7728 6 VGND
port 46 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 18548 20692
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/spm/runs/08-02_04-12/results/magic/spm.gds
string GDS_END 875588
string GDS_START 101976
<< end >>

